-- VideoBox.vhd

-- Generated using ACDS version 16.1 196

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity VideoBox is
	port (
		led_bus_export     : out   std_logic_vector(7 downto 0);                     --     led_bus.export
		memory_mem_a       : out   std_logic_vector(14 downto 0);                    --      memory.mem_a
		memory_mem_ba      : out   std_logic_vector(2 downto 0);                     --            .mem_ba
		memory_mem_ck      : out   std_logic;                                        --            .mem_ck
		memory_mem_ck_n    : out   std_logic;                                        --            .mem_ck_n
		memory_mem_cke     : out   std_logic;                                        --            .mem_cke
		memory_mem_cs_n    : out   std_logic;                                        --            .mem_cs_n
		memory_mem_ras_n   : out   std_logic;                                        --            .mem_ras_n
		memory_mem_cas_n   : out   std_logic;                                        --            .mem_cas_n
		memory_mem_we_n    : out   std_logic;                                        --            .mem_we_n
		memory_mem_reset_n : out   std_logic;                                        --            .mem_reset_n
		memory_mem_dq      : inout std_logic_vector(31 downto 0) := (others => '0'); --            .mem_dq
		memory_mem_dqs     : inout std_logic_vector(3 downto 0)  := (others => '0'); --            .mem_dqs
		memory_mem_dqs_n   : inout std_logic_vector(3 downto 0)  := (others => '0'); --            .mem_dqs_n
		memory_mem_odt     : out   std_logic;                                        --            .mem_odt
		memory_mem_dm      : out   std_logic_vector(3 downto 0);                     --            .mem_dm
		memory_oct_rzqin   : in    std_logic                     := '0';             --            .oct_rzqin
		ref_clock_clk      : in    std_logic                     := '0';             --   ref_clock.clk
		sdram_bus_addr     : out   std_logic_vector(12 downto 0);                    --   sdram_bus.addr
		sdram_bus_ba       : out   std_logic_vector(1 downto 0);                     --            .ba
		sdram_bus_cas_n    : out   std_logic;                                        --            .cas_n
		sdram_bus_cke      : out   std_logic;                                        --            .cke
		sdram_bus_cs_n     : out   std_logic;                                        --            .cs_n
		sdram_bus_dq       : inout std_logic_vector(15 downto 0) := (others => '0'); --            .dq
		sdram_bus_dqm      : out   std_logic_vector(1 downto 0);                     --            .dqm
		sdram_bus_ras_n    : out   std_logic;                                        --            .ras_n
		sdram_bus_we_n     : out   std_logic;                                        --            .we_n
		sdram_clock_clk    : out   std_logic;                                        -- sdram_clock.clk
		vga_bus_CLK        : out   std_logic;                                        --     vga_bus.CLK
		vga_bus_HS         : out   std_logic;                                        --            .HS
		vga_bus_VS         : out   std_logic;                                        --            .VS
		vga_bus_BLANK      : out   std_logic;                                        --            .BLANK
		vga_bus_SYNC       : out   std_logic;                                        --            .SYNC
		vga_bus_R          : out   std_logic_vector(7 downto 0);                     --            .R
		vga_bus_G          : out   std_logic_vector(7 downto 0);                     --            .G
		vga_bus_B          : out   std_logic_vector(7 downto 0)                      --            .B
	);
end entity VideoBox;

architecture rtl of VideoBox is
	component VideoBox_DMA_CONTROLLER_UPIS is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			stream_data          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			stream_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			stream_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			stream_valid         : in  std_logic                     := 'X';             -- valid
			stream_ready         : out std_logic;                                        -- ready
			slave_address        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			slave_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			slave_read           : in  std_logic                     := 'X';             -- read
			slave_write          : in  std_logic                     := 'X';             -- write
			slave_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_write         : out std_logic;                                        -- write
			master_writedata     : out std_logic_vector(15 downto 0)                     -- writedata
		);
	end component VideoBox_DMA_CONTROLLER_UPIS;

	component Image_Processing is
		port (
			avs_s0_address         : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			avs_s0_read            : in  std_logic                     := 'X';             -- read
			avs_s0_readdata        : out std_logic_vector(31 downto 0);                    -- readdata
			avs_s0_write           : in  std_logic                     := 'X';             -- write
			avs_s0_writedata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			asi_in0_data           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			asi_in0_ready          : out std_logic;                                        -- ready
			asi_in0_valid          : in  std_logic                     := 'X';             -- valid
			asi_in0_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			asi_in0_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			aso_out0_data          : out std_logic_vector(15 downto 0);                    -- data
			aso_out0_ready         : in  std_logic                     := 'X';             -- ready
			aso_out0_valid         : out std_logic;                                        -- valid
			aso_out0_endofpacket   : out std_logic;                                        -- endofpacket
			aso_out0_startofpacket : out std_logic;                                        -- startofpacket
			reset_reset            : in  std_logic                     := 'X';             -- reset
			clock_clk              : in  std_logic                     := 'X'              -- clk
		);
	end component Image_Processing;

	component Izbor_Prikaza_Slike is
		port (
			out_data               : out std_logic_vector(15 downto 0);                    -- data
			out_endofpacket        : out std_logic;                                        -- endofpacket
			out_ready              : in  std_logic                     := 'X';             -- ready
			out_startofpacket      : out std_logic;                                        -- startofpacket
			out_valid              : out std_logic;                                        -- valid
			in1_valid              : in  std_logic                     := 'X';             -- valid
			in1_startofpacket      : in  std_logic                     := 'X';             -- startofpacket
			in1_ready              : out std_logic;                                        -- ready
			in1_endofpacket        : in  std_logic                     := 'X';             -- endofpacket
			in1_data               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			in2_data               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			in2_ready              : out std_logic;                                        -- ready
			in2_valid              : in  std_logic                     := 'X';             -- valid
			in2_startofpacket      : in  std_logic                     := 'X';             -- startofpacket
			in2_endofpacket        : in  std_logic                     := 'X';             -- endofpacket
			clock_clk              : in  std_logic                     := 'X';             -- clk
			reset_reset            : in  std_logic                     := 'X';             -- reset
			izbor_slike_address    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			izbor_slike_write      : in  std_logic                     := 'X';             -- write
			izbor_slike_writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			izbor_slike_read       : in  std_logic                     := 'X';             -- read
			izbor_slike_readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			led_master_write       : out std_logic;                                        -- write
			led_master_writedata   : out std_logic_vector(7 downto 0);                     -- writedata
			led_master_waitrequest : in  std_logic                     := 'X'              -- waitrequest
		);
	end component Izbor_Prikaza_Slike;

	component Pozicioniranje_Piksela_u_SDRAM is
		port (
			reset_reset              : in  std_logic                     := 'X';             -- reset
			clock_clk                : in  std_logic                     := 'X';             -- clk
			out_piksel_data          : out std_logic_vector(15 downto 0);                    -- data
			out_piksel_endofpacket   : out std_logic;                                        -- endofpacket
			out_piksel_ready         : in  std_logic                     := 'X';             -- ready
			out_piksel_startofpacket : out std_logic;                                        -- startofpacket
			out_piksel_valid         : out std_logic;                                        -- valid
			in_piksel_ready          : out std_logic;                                        -- ready
			in_piksel_valid          : in  std_logic                     := 'X';             -- valid
			in_piksel_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			in_piksel_data           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			in_piksel_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_xy_valid              : in  std_logic                     := 'X';             -- valid
			in_xy_startofpacket      : in  std_logic                     := 'X';             -- startofpacket
			in_xy_endofpacket        : in  std_logic                     := 'X';             -- endofpacket
			in_xy_ready              : out std_logic;                                        -- ready
			in_xy_data               : in  std_logic_vector(31 downto 0) := (others => 'X')  -- data
		);
	end component Pozicioniranje_Piksela_u_SDRAM;

	component Transformacija_Slike is
		port (
			clock_clk              : in  std_logic                     := 'X';             -- clk
			reset_reset            : in  std_logic                     := 'X';             -- reset
			out_data               : out std_logic_vector(31 downto 0);                    -- data
			out_ready              : in  std_logic                     := 'X';             -- ready
			out_startofpacket      : out std_logic;                                        -- startofpacket
			out_endofpacket        : out std_logic;                                        -- endofpacket
			out_valid              : out std_logic;                                        -- valid
			avalon_slave_write     : in  std_logic                     := 'X';             -- write
			avalon_slave_writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			in_data                : in  std_logic_vector(63 downto 0) := (others => 'X'); -- data
			in_ready               : out std_logic;                                        -- ready
			in_startofpacket       : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket         : in  std_logic                     := 'X';             -- endofpacket
			in_valid               : in  std_logic                     := 'X'              -- valid
		);
	end component Transformacija_Slike;

	component VideoBox_affine_matrix is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			address     : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			address2    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk2        : in  std_logic                     := 'X';             -- clk
			reset2      : in  std_logic                     := 'X';             -- reset
			reset_req2  : in  std_logic                     := 'X';             -- reset_req
			freeze      : in  std_logic                     := 'X'              -- freeze
		);
	end component VideoBox_affine_matrix;

	component VideoBox_dma_afina_matrica_citanje is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_arbiterlock   : out std_logic;                                        -- lock
			master_read          : out std_logic;                                        -- read
			master_readdata      : in  std_logic_vector(63 downto 0) := (others => 'X'); -- readdata
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			slave_address        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			slave_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			slave_read           : in  std_logic                     := 'X';             -- read
			slave_write          : in  std_logic                     := 'X';             -- write
			slave_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			stream_ready         : in  std_logic                     := 'X';             -- ready
			stream_data          : out std_logic_vector(63 downto 0);                    -- data
			stream_startofpacket : out std_logic;                                        -- startofpacket
			stream_endofpacket   : out std_logic;                                        -- endofpacket
			stream_valid         : out std_logic                                         -- valid
		);
	end component VideoBox_dma_afina_matrica_citanje;

	component VideoBox_hps is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			mem_a          : out   std_logic_vector(14 downto 0);                    -- mem_a
			mem_ba         : out   std_logic_vector(2 downto 0);                     -- mem_ba
			mem_ck         : out   std_logic;                                        -- mem_ck
			mem_ck_n       : out   std_logic;                                        -- mem_ck_n
			mem_cke        : out   std_logic;                                        -- mem_cke
			mem_cs_n       : out   std_logic;                                        -- mem_cs_n
			mem_ras_n      : out   std_logic;                                        -- mem_ras_n
			mem_cas_n      : out   std_logic;                                        -- mem_cas_n
			mem_we_n       : out   std_logic;                                        -- mem_we_n
			mem_reset_n    : out   std_logic;                                        -- mem_reset_n
			mem_dq         : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs        : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n      : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
			mem_odt        : out   std_logic;                                        -- mem_odt
			mem_dm         : out   std_logic_vector(3 downto 0);                     -- mem_dm
			oct_rzqin      : in    std_logic                     := 'X';             -- oct_rzqin
			h2f_rst_n      : out   std_logic;                                        -- reset_n
			h2f_axi_clk    : in    std_logic                     := 'X';             -- clk
			h2f_AWID       : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_AWADDR     : out   std_logic_vector(29 downto 0);                    -- awaddr
			h2f_AWLEN      : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_AWSIZE     : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_AWBURST    : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_AWLOCK     : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_AWCACHE    : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_AWPROT     : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_AWVALID    : out   std_logic;                                        -- awvalid
			h2f_AWREADY    : in    std_logic                     := 'X';             -- awready
			h2f_WID        : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_WDATA      : out   std_logic_vector(63 downto 0);                    -- wdata
			h2f_WSTRB      : out   std_logic_vector(7 downto 0);                     -- wstrb
			h2f_WLAST      : out   std_logic;                                        -- wlast
			h2f_WVALID     : out   std_logic;                                        -- wvalid
			h2f_WREADY     : in    std_logic                     := 'X';             -- wready
			h2f_BID        : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_BRESP      : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_BVALID     : in    std_logic                     := 'X';             -- bvalid
			h2f_BREADY     : out   std_logic;                                        -- bready
			h2f_ARID       : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_ARADDR     : out   std_logic_vector(29 downto 0);                    -- araddr
			h2f_ARLEN      : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_ARSIZE     : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_ARBURST    : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_ARLOCK     : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_ARCACHE    : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_ARPROT     : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_ARVALID    : out   std_logic;                                        -- arvalid
			h2f_ARREADY    : in    std_logic                     := 'X';             -- arready
			h2f_RID        : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_RDATA      : in    std_logic_vector(63 downto 0) := (others => 'X'); -- rdata
			h2f_RRESP      : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_RLAST      : in    std_logic                     := 'X';             -- rlast
			h2f_RVALID     : in    std_logic                     := 'X';             -- rvalid
			h2f_RREADY     : out   std_logic;                                        -- rready
			h2f_lw_axi_clk : in    std_logic                     := 'X';             -- clk
			h2f_lw_AWID    : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_lw_AWADDR  : out   std_logic_vector(20 downto 0);                    -- awaddr
			h2f_lw_AWLEN   : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_lw_AWSIZE  : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_lw_AWBURST : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_lw_AWLOCK  : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_lw_AWCACHE : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_lw_AWPROT  : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_lw_AWVALID : out   std_logic;                                        -- awvalid
			h2f_lw_AWREADY : in    std_logic                     := 'X';             -- awready
			h2f_lw_WID     : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_lw_WDATA   : out   std_logic_vector(31 downto 0);                    -- wdata
			h2f_lw_WSTRB   : out   std_logic_vector(3 downto 0);                     -- wstrb
			h2f_lw_WLAST   : out   std_logic;                                        -- wlast
			h2f_lw_WVALID  : out   std_logic;                                        -- wvalid
			h2f_lw_WREADY  : in    std_logic                     := 'X';             -- wready
			h2f_lw_BID     : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_lw_BRESP   : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_lw_BVALID  : in    std_logic                     := 'X';             -- bvalid
			h2f_lw_BREADY  : out   std_logic;                                        -- bready
			h2f_lw_ARID    : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_lw_ARADDR  : out   std_logic_vector(20 downto 0);                    -- araddr
			h2f_lw_ARLEN   : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_lw_ARSIZE  : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_lw_ARBURST : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_lw_ARLOCK  : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_lw_ARCACHE : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_lw_ARPROT  : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_lw_ARVALID : out   std_logic;                                        -- arvalid
			h2f_lw_ARREADY : in    std_logic                     := 'X';             -- arready
			h2f_lw_RID     : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_lw_RDATA   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			h2f_lw_RRESP   : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_lw_RLAST   : in    std_logic                     := 'X';             -- rlast
			h2f_lw_RVALID  : in    std_logic                     := 'X';             -- rvalid
			h2f_lw_RREADY  : out   std_logic                                         -- rready
		);
	end component VideoBox_hps;

	component VideoBox_led_indication_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component VideoBox_led_indication_0;

	component VideoBox_sdram_controller is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component VideoBox_sdram_controller;

	component VideoBox_sys_sdram_pll is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			sys_clk_clk        : out std_logic;        -- clk
			sdram_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component VideoBox_sys_sdram_pll;

	component VideoBox_vga_pll is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component VideoBox_vga_pll;

	component VideoBox_vide_dma_controller is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_arbiterlock   : out std_logic;                                        -- lock
			master_read          : out std_logic;                                        -- read
			master_readdata      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			slave_address        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			slave_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			slave_read           : in  std_logic                     := 'X';             -- read
			slave_write          : in  std_logic                     := 'X';             -- write
			slave_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			stream_ready         : in  std_logic                     := 'X';             -- ready
			stream_data          : out std_logic_vector(15 downto 0);                    -- data
			stream_startofpacket : out std_logic;                                        -- startofpacket
			stream_endofpacket   : out std_logic;                                        -- endofpacket
			stream_valid         : out std_logic                                         -- valid
		);
	end component VideoBox_vide_dma_controller;

	component VideoBox_vide_dma_controller_CITANJE is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_arbiterlock   : out std_logic;                                        -- lock
			master_read          : out std_logic;                                        -- read
			master_readdata      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			slave_address        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			slave_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			slave_read           : in  std_logic                     := 'X';             -- read
			slave_write          : in  std_logic                     := 'X';             -- write
			slave_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			stream_ready         : in  std_logic                     := 'X';             -- ready
			stream_data          : out std_logic_vector(15 downto 0);                    -- data
			stream_startofpacket : out std_logic;                                        -- startofpacket
			stream_endofpacket   : out std_logic;                                        -- endofpacket
			stream_valid         : out std_logic                                         -- valid
		);
	end component VideoBox_vide_dma_controller_CITANJE;

	component VideoBox_video_dual_clock_buffer is
		port (
			clk_stream_in            : in  std_logic                     := 'X';             -- clk
			reset_stream_in          : in  std_logic                     := 'X';             -- reset
			clk_stream_out           : in  std_logic                     := 'X';             -- clk
			reset_stream_out         : in  std_logic                     := 'X';             -- reset
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_data           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(15 downto 0)                     -- data
		);
	end component VideoBox_video_dual_clock_buffer;

	component VideoBox_video_rgb_resampler_0 is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_data           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(29 downto 0)                     -- data
		);
	end component VideoBox_video_rgb_resampler_0;

	component VideoBox_video_vga_controller is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			data          : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			startofpacket : in  std_logic                     := 'X';             -- startofpacket
			endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			valid         : in  std_logic                     := 'X';             -- valid
			ready         : out std_logic;                                        -- ready
			VGA_CLK       : out std_logic;                                        -- export
			VGA_HS        : out std_logic;                                        -- export
			VGA_VS        : out std_logic;                                        -- export
			VGA_BLANK     : out std_logic;                                        -- export
			VGA_SYNC      : out std_logic;                                        -- export
			VGA_R         : out std_logic_vector(7 downto 0);                     -- export
			VGA_G         : out std_logic_vector(7 downto 0);                     -- export
			VGA_B         : out std_logic_vector(7 downto 0)                      -- export
		);
	end component VideoBox_video_vga_controller;

	component VideoBox_mm_interconnect_0 is
		port (
			hps_h2f_axi_master_awid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			hps_h2f_axi_master_awaddr                                      : in  std_logic_vector(29 downto 0) := (others => 'X'); -- awaddr
			hps_h2f_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			hps_h2f_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			hps_h2f_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			hps_h2f_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			hps_h2f_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			hps_h2f_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			hps_h2f_axi_master_awvalid                                     : in  std_logic                     := 'X';             -- awvalid
			hps_h2f_axi_master_awready                                     : out std_logic;                                        -- awready
			hps_h2f_axi_master_wid                                         : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			hps_h2f_axi_master_wdata                                       : in  std_logic_vector(63 downto 0) := (others => 'X'); -- wdata
			hps_h2f_axi_master_wstrb                                       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wstrb
			hps_h2f_axi_master_wlast                                       : in  std_logic                     := 'X';             -- wlast
			hps_h2f_axi_master_wvalid                                      : in  std_logic                     := 'X';             -- wvalid
			hps_h2f_axi_master_wready                                      : out std_logic;                                        -- wready
			hps_h2f_axi_master_bid                                         : out std_logic_vector(11 downto 0);                    -- bid
			hps_h2f_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                     -- bresp
			hps_h2f_axi_master_bvalid                                      : out std_logic;                                        -- bvalid
			hps_h2f_axi_master_bready                                      : in  std_logic                     := 'X';             -- bready
			hps_h2f_axi_master_arid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			hps_h2f_axi_master_araddr                                      : in  std_logic_vector(29 downto 0) := (others => 'X'); -- araddr
			hps_h2f_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			hps_h2f_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			hps_h2f_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			hps_h2f_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			hps_h2f_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			hps_h2f_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			hps_h2f_axi_master_arvalid                                     : in  std_logic                     := 'X';             -- arvalid
			hps_h2f_axi_master_arready                                     : out std_logic;                                        -- arready
			hps_h2f_axi_master_rid                                         : out std_logic_vector(11 downto 0);                    -- rid
			hps_h2f_axi_master_rdata                                       : out std_logic_vector(63 downto 0);                    -- rdata
			hps_h2f_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                     -- rresp
			hps_h2f_axi_master_rlast                                       : out std_logic;                                        -- rlast
			hps_h2f_axi_master_rvalid                                      : out std_logic;                                        -- rvalid
			hps_h2f_axi_master_rready                                      : in  std_logic                     := 'X';             -- rready
			sys_sdram_pll_sys_clk_clk                                      : in  std_logic                     := 'X';             -- clk
			hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			vide_dma_controller_reset_reset_bridge_in_reset_reset          : in  std_logic                     := 'X';             -- reset
			dma_afina_matrica_citanje_avalon_dma_master_address            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			dma_afina_matrica_citanje_avalon_dma_master_waitrequest        : out std_logic;                                        -- waitrequest
			dma_afina_matrica_citanje_avalon_dma_master_read               : in  std_logic                     := 'X';             -- read
			dma_afina_matrica_citanje_avalon_dma_master_readdata           : out std_logic_vector(63 downto 0);                    -- readdata
			dma_afina_matrica_citanje_avalon_dma_master_readdatavalid      : out std_logic;                                        -- readdatavalid
			dma_afina_matrica_citanje_avalon_dma_master_lock               : in  std_logic                     := 'X';             -- lock
			DMA_CONTROLLER_UPIS_avalon_dma_master_address                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			DMA_CONTROLLER_UPIS_avalon_dma_master_waitrequest              : out std_logic;                                        -- waitrequest
			DMA_CONTROLLER_UPIS_avalon_dma_master_write                    : in  std_logic                     := 'X';             -- write
			DMA_CONTROLLER_UPIS_avalon_dma_master_writedata                : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			vide_dma_controller_avalon_dma_master_address                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			vide_dma_controller_avalon_dma_master_waitrequest              : out std_logic;                                        -- waitrequest
			vide_dma_controller_avalon_dma_master_read                     : in  std_logic                     := 'X';             -- read
			vide_dma_controller_avalon_dma_master_readdata                 : out std_logic_vector(15 downto 0);                    -- readdata
			vide_dma_controller_avalon_dma_master_readdatavalid            : out std_logic;                                        -- readdatavalid
			vide_dma_controller_avalon_dma_master_lock                     : in  std_logic                     := 'X';             -- lock
			vide_dma_controller_CITANJE_avalon_dma_master_address          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			vide_dma_controller_CITANJE_avalon_dma_master_waitrequest      : out std_logic;                                        -- waitrequest
			vide_dma_controller_CITANJE_avalon_dma_master_read             : in  std_logic                     := 'X';             -- read
			vide_dma_controller_CITANJE_avalon_dma_master_readdata         : out std_logic_vector(15 downto 0);                    -- readdata
			vide_dma_controller_CITANJE_avalon_dma_master_readdatavalid    : out std_logic;                                        -- readdatavalid
			vide_dma_controller_CITANJE_avalon_dma_master_lock             : in  std_logic                     := 'X';             -- lock
			vide_dma_controller_CITANJE_0_avalon_dma_master_address        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			vide_dma_controller_CITANJE_0_avalon_dma_master_waitrequest    : out std_logic;                                        -- waitrequest
			vide_dma_controller_CITANJE_0_avalon_dma_master_read           : in  std_logic                     := 'X';             -- read
			vide_dma_controller_CITANJE_0_avalon_dma_master_readdata       : out std_logic_vector(15 downto 0);                    -- readdata
			vide_dma_controller_CITANJE_0_avalon_dma_master_readdatavalid  : out std_logic;                                        -- readdatavalid
			vide_dma_controller_CITANJE_0_avalon_dma_master_lock           : in  std_logic                     := 'X';             -- lock
			affine_matrix_s1_address                                       : out std_logic_vector(9 downto 0);                     -- address
			affine_matrix_s1_write                                         : out std_logic;                                        -- write
			affine_matrix_s1_readdata                                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			affine_matrix_s1_writedata                                     : out std_logic_vector(31 downto 0);                    -- writedata
			affine_matrix_s1_byteenable                                    : out std_logic_vector(3 downto 0);                     -- byteenable
			affine_matrix_s1_chipselect                                    : out std_logic;                                        -- chipselect
			affine_matrix_s1_clken                                         : out std_logic;                                        -- clken
			sdram_controller_s1_address                                    : out std_logic_vector(24 downto 0);                    -- address
			sdram_controller_s1_write                                      : out std_logic;                                        -- write
			sdram_controller_s1_read                                       : out std_logic;                                        -- read
			sdram_controller_s1_readdata                                   : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_controller_s1_writedata                                  : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_controller_s1_byteenable                                 : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_controller_s1_readdatavalid                              : in  std_logic                     := 'X';             -- readdatavalid
			sdram_controller_s1_waitrequest                                : in  std_logic                     := 'X';             -- waitrequest
			sdram_controller_s1_chipselect                                 : out std_logic                                         -- chipselect
		);
	end component VideoBox_mm_interconnect_0;

	component VideoBox_mm_interconnect_1 is
		port (
			hps_h2f_lw_axi_master_awid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			hps_h2f_lw_axi_master_awaddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- awaddr
			hps_h2f_lw_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			hps_h2f_lw_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			hps_h2f_lw_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			hps_h2f_lw_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			hps_h2f_lw_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			hps_h2f_lw_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			hps_h2f_lw_axi_master_awvalid                                     : in  std_logic                     := 'X';             -- awvalid
			hps_h2f_lw_axi_master_awready                                     : out std_logic;                                        -- awready
			hps_h2f_lw_axi_master_wid                                         : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			hps_h2f_lw_axi_master_wdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			hps_h2f_lw_axi_master_wstrb                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			hps_h2f_lw_axi_master_wlast                                       : in  std_logic                     := 'X';             -- wlast
			hps_h2f_lw_axi_master_wvalid                                      : in  std_logic                     := 'X';             -- wvalid
			hps_h2f_lw_axi_master_wready                                      : out std_logic;                                        -- wready
			hps_h2f_lw_axi_master_bid                                         : out std_logic_vector(11 downto 0);                    -- bid
			hps_h2f_lw_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                     -- bresp
			hps_h2f_lw_axi_master_bvalid                                      : out std_logic;                                        -- bvalid
			hps_h2f_lw_axi_master_bready                                      : in  std_logic                     := 'X';             -- bready
			hps_h2f_lw_axi_master_arid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			hps_h2f_lw_axi_master_araddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- araddr
			hps_h2f_lw_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			hps_h2f_lw_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			hps_h2f_lw_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			hps_h2f_lw_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			hps_h2f_lw_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			hps_h2f_lw_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			hps_h2f_lw_axi_master_arvalid                                     : in  std_logic                     := 'X';             -- arvalid
			hps_h2f_lw_axi_master_arready                                     : out std_logic;                                        -- arready
			hps_h2f_lw_axi_master_rid                                         : out std_logic_vector(11 downto 0);                    -- rid
			hps_h2f_lw_axi_master_rdata                                       : out std_logic_vector(31 downto 0);                    -- rdata
			hps_h2f_lw_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                     -- rresp
			hps_h2f_lw_axi_master_rlast                                       : out std_logic;                                        -- rlast
			hps_h2f_lw_axi_master_rvalid                                      : out std_logic;                                        -- rvalid
			hps_h2f_lw_axi_master_rready                                      : in  std_logic                     := 'X';             -- rready
			sys_sdram_pll_sys_clk_clk                                         : in  std_logic                     := 'X';             -- clk
			hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			vide_dma_controller_reset_reset_bridge_in_reset_reset             : in  std_logic                     := 'X';             -- reset
			DMA_CONTROLLER_UPIS_avalon_dma_control_slave_address              : out std_logic_vector(1 downto 0);                     -- address
			DMA_CONTROLLER_UPIS_avalon_dma_control_slave_write                : out std_logic;                                        -- write
			DMA_CONTROLLER_UPIS_avalon_dma_control_slave_read                 : out std_logic;                                        -- read
			DMA_CONTROLLER_UPIS_avalon_dma_control_slave_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			DMA_CONTROLLER_UPIS_avalon_dma_control_slave_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			DMA_CONTROLLER_UPIS_avalon_dma_control_slave_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			Image_Processing_0_s0_address                                     : out std_logic_vector(7 downto 0);                     -- address
			Image_Processing_0_s0_write                                       : out std_logic;                                        -- write
			Image_Processing_0_s0_read                                        : out std_logic;                                        -- read
			Image_Processing_0_s0_readdata                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Image_Processing_0_s0_writedata                                   : out std_logic_vector(31 downto 0);                    -- writedata
			Izbor_Prikaza_Slike_0_izbor_slike_address                         : out std_logic_vector(7 downto 0);                     -- address
			Izbor_Prikaza_Slike_0_izbor_slike_write                           : out std_logic;                                        -- write
			Izbor_Prikaza_Slike_0_izbor_slike_read                            : out std_logic;                                        -- read
			Izbor_Prikaza_Slike_0_izbor_slike_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Izbor_Prikaza_Slike_0_izbor_slike_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			vide_dma_controller_avalon_dma_control_slave_address              : out std_logic_vector(1 downto 0);                     -- address
			vide_dma_controller_avalon_dma_control_slave_write                : out std_logic;                                        -- write
			vide_dma_controller_avalon_dma_control_slave_read                 : out std_logic;                                        -- read
			vide_dma_controller_avalon_dma_control_slave_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			vide_dma_controller_avalon_dma_control_slave_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			vide_dma_controller_avalon_dma_control_slave_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			vide_dma_controller_CITANJE_avalon_dma_control_slave_address      : out std_logic_vector(1 downto 0);                     -- address
			vide_dma_controller_CITANJE_avalon_dma_control_slave_write        : out std_logic;                                        -- write
			vide_dma_controller_CITANJE_avalon_dma_control_slave_read         : out std_logic;                                        -- read
			vide_dma_controller_CITANJE_avalon_dma_control_slave_readdata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			vide_dma_controller_CITANJE_avalon_dma_control_slave_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			vide_dma_controller_CITANJE_avalon_dma_control_slave_byteenable   : out std_logic_vector(3 downto 0);                     -- byteenable
			vide_dma_controller_CITANJE_0_avalon_dma_control_slave_address    : out std_logic_vector(1 downto 0);                     -- address
			vide_dma_controller_CITANJE_0_avalon_dma_control_slave_write      : out std_logic;                                        -- write
			vide_dma_controller_CITANJE_0_avalon_dma_control_slave_read       : out std_logic;                                        -- read
			vide_dma_controller_CITANJE_0_avalon_dma_control_slave_readdata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			vide_dma_controller_CITANJE_0_avalon_dma_control_slave_writedata  : out std_logic_vector(31 downto 0);                    -- writedata
			vide_dma_controller_CITANJE_0_avalon_dma_control_slave_byteenable : out std_logic_vector(3 downto 0)                      -- byteenable
		);
	end component VideoBox_mm_interconnect_1;

	component VideoBox_mm_interconnect_2 is
		port (
			sys_sdram_pll_sys_clk_clk                               : in  std_logic                     := 'X';             -- clk
			Izbor_Prikaza_Slike_0_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			Izbor_Prikaza_Slike_0_led_master_waitrequest            : out std_logic;                                        -- waitrequest
			Izbor_Prikaza_Slike_0_led_master_write                  : in  std_logic                     := 'X';             -- write
			Izbor_Prikaza_Slike_0_led_master_writedata              : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			led_indication_0_s1_address                             : out std_logic_vector(1 downto 0);                     -- address
			led_indication_0_s1_write                               : out std_logic;                                        -- write
			led_indication_0_s1_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_indication_0_s1_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			led_indication_0_s1_chipselect                          : out std_logic                                         -- chipselect
		);
	end component VideoBox_mm_interconnect_2;

	component videobox_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component videobox_rst_controller;

	component videobox_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component videobox_rst_controller_001;

	signal video_dual_clock_buffer_avalon_dc_buffer_source_valid                               : std_logic;                     -- video_dual_clock_buffer:stream_out_valid -> video_rgb_resampler_0:stream_in_valid
	signal video_dual_clock_buffer_avalon_dc_buffer_source_data                                : std_logic_vector(15 downto 0); -- video_dual_clock_buffer:stream_out_data -> video_rgb_resampler_0:stream_in_data
	signal video_dual_clock_buffer_avalon_dc_buffer_source_ready                               : std_logic;                     -- video_rgb_resampler_0:stream_in_ready -> video_dual_clock_buffer:stream_out_ready
	signal video_dual_clock_buffer_avalon_dc_buffer_source_startofpacket                       : std_logic;                     -- video_dual_clock_buffer:stream_out_startofpacket -> video_rgb_resampler_0:stream_in_startofpacket
	signal video_dual_clock_buffer_avalon_dc_buffer_source_endofpacket                         : std_logic;                     -- video_dual_clock_buffer:stream_out_endofpacket -> video_rgb_resampler_0:stream_in_endofpacket
	signal vide_dma_controller_citanje_0_avalon_pixel_source_valid                             : std_logic;                     -- vide_dma_controller_CITANJE_0:stream_valid -> Image_Processing_0:asi_in0_valid
	signal vide_dma_controller_citanje_0_avalon_pixel_source_data                              : std_logic_vector(15 downto 0); -- vide_dma_controller_CITANJE_0:stream_data -> Image_Processing_0:asi_in0_data
	signal vide_dma_controller_citanje_0_avalon_pixel_source_ready                             : std_logic;                     -- Image_Processing_0:asi_in0_ready -> vide_dma_controller_CITANJE_0:stream_ready
	signal vide_dma_controller_citanje_0_avalon_pixel_source_startofpacket                     : std_logic;                     -- vide_dma_controller_CITANJE_0:stream_startofpacket -> Image_Processing_0:asi_in0_startofpacket
	signal vide_dma_controller_citanje_0_avalon_pixel_source_endofpacket                       : std_logic;                     -- vide_dma_controller_CITANJE_0:stream_endofpacket -> Image_Processing_0:asi_in0_endofpacket
	signal vide_dma_controller_citanje_avalon_pixel_source_valid                               : std_logic;                     -- vide_dma_controller_CITANJE:stream_valid -> Izbor_Prikaza_Slike_0:in1_valid
	signal vide_dma_controller_citanje_avalon_pixel_source_data                                : std_logic_vector(15 downto 0); -- vide_dma_controller_CITANJE:stream_data -> Izbor_Prikaza_Slike_0:in1_data
	signal vide_dma_controller_citanje_avalon_pixel_source_ready                               : std_logic;                     -- Izbor_Prikaza_Slike_0:in1_ready -> vide_dma_controller_CITANJE:stream_ready
	signal vide_dma_controller_citanje_avalon_pixel_source_startofpacket                       : std_logic;                     -- vide_dma_controller_CITANJE:stream_startofpacket -> Izbor_Prikaza_Slike_0:in1_startofpacket
	signal vide_dma_controller_citanje_avalon_pixel_source_endofpacket                         : std_logic;                     -- vide_dma_controller_CITANJE:stream_endofpacket -> Izbor_Prikaza_Slike_0:in1_endofpacket
	signal vide_dma_controller_avalon_pixel_source_valid                                       : std_logic;                     -- vide_dma_controller:stream_valid -> Izbor_Prikaza_Slike_0:in2_valid
	signal vide_dma_controller_avalon_pixel_source_data                                        : std_logic_vector(15 downto 0); -- vide_dma_controller:stream_data -> Izbor_Prikaza_Slike_0:in2_data
	signal vide_dma_controller_avalon_pixel_source_ready                                       : std_logic;                     -- Izbor_Prikaza_Slike_0:in2_ready -> vide_dma_controller:stream_ready
	signal vide_dma_controller_avalon_pixel_source_startofpacket                               : std_logic;                     -- vide_dma_controller:stream_startofpacket -> Izbor_Prikaza_Slike_0:in2_startofpacket
	signal vide_dma_controller_avalon_pixel_source_endofpacket                                 : std_logic;                     -- vide_dma_controller:stream_endofpacket -> Izbor_Prikaza_Slike_0:in2_endofpacket
	signal dma_afina_matrica_citanje_avalon_pixel_source_valid                                 : std_logic;                     -- dma_afina_matrica_citanje:stream_valid -> Transformacija_Pozicije_Piksela:in_valid
	signal dma_afina_matrica_citanje_avalon_pixel_source_data                                  : std_logic_vector(63 downto 0); -- dma_afina_matrica_citanje:stream_data -> Transformacija_Pozicije_Piksela:in_data
	signal dma_afina_matrica_citanje_avalon_pixel_source_ready                                 : std_logic;                     -- Transformacija_Pozicije_Piksela:in_ready -> dma_afina_matrica_citanje:stream_ready
	signal dma_afina_matrica_citanje_avalon_pixel_source_startofpacket                         : std_logic;                     -- dma_afina_matrica_citanje:stream_startofpacket -> Transformacija_Pozicije_Piksela:in_startofpacket
	signal dma_afina_matrica_citanje_avalon_pixel_source_endofpacket                           : std_logic;                     -- dma_afina_matrica_citanje:stream_endofpacket -> Transformacija_Pozicije_Piksela:in_endofpacket
	signal video_rgb_resampler_0_avalon_rgb_source_valid                                       : std_logic;                     -- video_rgb_resampler_0:stream_out_valid -> video_vga_controller:valid
	signal video_rgb_resampler_0_avalon_rgb_source_data                                        : std_logic_vector(29 downto 0); -- video_rgb_resampler_0:stream_out_data -> video_vga_controller:data
	signal video_rgb_resampler_0_avalon_rgb_source_ready                                       : std_logic;                     -- video_vga_controller:ready -> video_rgb_resampler_0:stream_out_ready
	signal video_rgb_resampler_0_avalon_rgb_source_startofpacket                               : std_logic;                     -- video_rgb_resampler_0:stream_out_startofpacket -> video_vga_controller:startofpacket
	signal video_rgb_resampler_0_avalon_rgb_source_endofpacket                                 : std_logic;                     -- video_rgb_resampler_0:stream_out_endofpacket -> video_vga_controller:endofpacket
	signal izbor_prikaza_slike_0_out_valid                                                     : std_logic;                     -- Izbor_Prikaza_Slike_0:out_valid -> video_dual_clock_buffer:stream_in_valid
	signal izbor_prikaza_slike_0_out_data                                                      : std_logic_vector(15 downto 0); -- Izbor_Prikaza_Slike_0:out_data -> video_dual_clock_buffer:stream_in_data
	signal izbor_prikaza_slike_0_out_ready                                                     : std_logic;                     -- video_dual_clock_buffer:stream_in_ready -> Izbor_Prikaza_Slike_0:out_ready
	signal izbor_prikaza_slike_0_out_startofpacket                                             : std_logic;                     -- Izbor_Prikaza_Slike_0:out_startofpacket -> video_dual_clock_buffer:stream_in_startofpacket
	signal izbor_prikaza_slike_0_out_endofpacket                                               : std_logic;                     -- Izbor_Prikaza_Slike_0:out_endofpacket -> video_dual_clock_buffer:stream_in_endofpacket
	signal image_processing_0_out0_valid                                                       : std_logic;                     -- Image_Processing_0:aso_out0_valid -> DMA_CONTROLLER_UPIS:stream_valid
	signal image_processing_0_out0_data                                                        : std_logic_vector(15 downto 0); -- Image_Processing_0:aso_out0_data -> DMA_CONTROLLER_UPIS:stream_data
	signal image_processing_0_out0_ready                                                       : std_logic;                     -- DMA_CONTROLLER_UPIS:stream_ready -> Image_Processing_0:aso_out0_ready
	signal image_processing_0_out0_startofpacket                                               : std_logic;                     -- Image_Processing_0:aso_out0_startofpacket -> DMA_CONTROLLER_UPIS:stream_startofpacket
	signal image_processing_0_out0_endofpacket                                                 : std_logic;                     -- Image_Processing_0:aso_out0_endofpacket -> DMA_CONTROLLER_UPIS:stream_endofpacket
	signal transformacija_pozicije_piksela_xy_out_valid                                        : std_logic;                     -- Transformacija_Pozicije_Piksela:out_valid -> Pozicioniranje_Piksela_u_SDRAM_0:in_xy_valid
	signal transformacija_pozicije_piksela_xy_out_data                                         : std_logic_vector(31 downto 0); -- Transformacija_Pozicije_Piksela:out_data -> Pozicioniranje_Piksela_u_SDRAM_0:in_xy_data
	signal transformacija_pozicije_piksela_xy_out_ready                                        : std_logic;                     -- Pozicioniranje_Piksela_u_SDRAM_0:in_xy_ready -> Transformacija_Pozicije_Piksela:out_ready
	signal transformacija_pozicije_piksela_xy_out_startofpacket                                : std_logic;                     -- Transformacija_Pozicije_Piksela:out_startofpacket -> Pozicioniranje_Piksela_u_SDRAM_0:in_xy_startofpacket
	signal transformacija_pozicije_piksela_xy_out_endofpacket                                  : std_logic;                     -- Transformacija_Pozicije_Piksela:out_endofpacket -> Pozicioniranje_Piksela_u_SDRAM_0:in_xy_endofpacket
	signal vga_pll_outclk0_clk                                                                 : std_logic;                     -- vga_pll:outclk_0 -> [rst_controller_001:clk, video_dual_clock_buffer:clk_stream_out, video_rgb_resampler_0:clk, video_vga_controller:clk]
	signal sys_sdram_pll_sys_clk_clk                                                           : std_logic;                     -- sys_sdram_pll:sys_clk_clk -> [DMA_CONTROLLER_UPIS:clk, Image_Processing_0:clock_clk, Izbor_Prikaza_Slike_0:clock_clk, Pozicioniranje_Piksela_u_SDRAM_0:clock_clk, Transformacija_Pozicije_Piksela:clock_clk, affine_matrix:clk, affine_matrix:clk2, dma_afina_matrica_citanje:clk, hps:h2f_axi_clk, hps:h2f_lw_axi_clk, led_indication_0:clk, mm_interconnect_0:sys_sdram_pll_sys_clk_clk, mm_interconnect_1:sys_sdram_pll_sys_clk_clk, mm_interconnect_2:sys_sdram_pll_sys_clk_clk, rst_controller:clk, rst_controller_002:clk, sdram_controller:clk, vga_pll:refclk, vide_dma_controller:clk, vide_dma_controller_CITANJE:clk, vide_dma_controller_CITANJE_0:clk, video_dual_clock_buffer:clk_stream_in]
	signal hps_h2f_reset_reset                                                                 : std_logic;                     -- hps:h2f_rst_n -> hps_h2f_reset_reset:in
	signal sys_sdram_pll_reset_source_reset                                                    : std_logic;                     -- sys_sdram_pll:reset_source_reset -> [rst_controller:reset_in0, rst_controller_001:reset_in0, vga_pll:rst]
	signal vide_dma_controller_avalon_dma_master_waitrequest                                   : std_logic;                     -- mm_interconnect_0:vide_dma_controller_avalon_dma_master_waitrequest -> vide_dma_controller:master_waitrequest
	signal vide_dma_controller_avalon_dma_master_readdata                                      : std_logic_vector(15 downto 0); -- mm_interconnect_0:vide_dma_controller_avalon_dma_master_readdata -> vide_dma_controller:master_readdata
	signal vide_dma_controller_avalon_dma_master_address                                       : std_logic_vector(31 downto 0); -- vide_dma_controller:master_address -> mm_interconnect_0:vide_dma_controller_avalon_dma_master_address
	signal vide_dma_controller_avalon_dma_master_read                                          : std_logic;                     -- vide_dma_controller:master_read -> mm_interconnect_0:vide_dma_controller_avalon_dma_master_read
	signal vide_dma_controller_avalon_dma_master_readdatavalid                                 : std_logic;                     -- mm_interconnect_0:vide_dma_controller_avalon_dma_master_readdatavalid -> vide_dma_controller:master_readdatavalid
	signal vide_dma_controller_avalon_dma_master_lock                                          : std_logic;                     -- vide_dma_controller:master_arbiterlock -> mm_interconnect_0:vide_dma_controller_avalon_dma_master_lock
	signal vide_dma_controller_citanje_avalon_dma_master_waitrequest                           : std_logic;                     -- mm_interconnect_0:vide_dma_controller_CITANJE_avalon_dma_master_waitrequest -> vide_dma_controller_CITANJE:master_waitrequest
	signal vide_dma_controller_citanje_avalon_dma_master_readdata                              : std_logic_vector(15 downto 0); -- mm_interconnect_0:vide_dma_controller_CITANJE_avalon_dma_master_readdata -> vide_dma_controller_CITANJE:master_readdata
	signal vide_dma_controller_citanje_avalon_dma_master_address                               : std_logic_vector(31 downto 0); -- vide_dma_controller_CITANJE:master_address -> mm_interconnect_0:vide_dma_controller_CITANJE_avalon_dma_master_address
	signal vide_dma_controller_citanje_avalon_dma_master_read                                  : std_logic;                     -- vide_dma_controller_CITANJE:master_read -> mm_interconnect_0:vide_dma_controller_CITANJE_avalon_dma_master_read
	signal vide_dma_controller_citanje_avalon_dma_master_readdatavalid                         : std_logic;                     -- mm_interconnect_0:vide_dma_controller_CITANJE_avalon_dma_master_readdatavalid -> vide_dma_controller_CITANJE:master_readdatavalid
	signal vide_dma_controller_citanje_avalon_dma_master_lock                                  : std_logic;                     -- vide_dma_controller_CITANJE:master_arbiterlock -> mm_interconnect_0:vide_dma_controller_CITANJE_avalon_dma_master_lock
	signal vide_dma_controller_citanje_0_avalon_dma_master_waitrequest                         : std_logic;                     -- mm_interconnect_0:vide_dma_controller_CITANJE_0_avalon_dma_master_waitrequest -> vide_dma_controller_CITANJE_0:master_waitrequest
	signal vide_dma_controller_citanje_0_avalon_dma_master_readdata                            : std_logic_vector(15 downto 0); -- mm_interconnect_0:vide_dma_controller_CITANJE_0_avalon_dma_master_readdata -> vide_dma_controller_CITANJE_0:master_readdata
	signal vide_dma_controller_citanje_0_avalon_dma_master_address                             : std_logic_vector(31 downto 0); -- vide_dma_controller_CITANJE_0:master_address -> mm_interconnect_0:vide_dma_controller_CITANJE_0_avalon_dma_master_address
	signal vide_dma_controller_citanje_0_avalon_dma_master_read                                : std_logic;                     -- vide_dma_controller_CITANJE_0:master_read -> mm_interconnect_0:vide_dma_controller_CITANJE_0_avalon_dma_master_read
	signal vide_dma_controller_citanje_0_avalon_dma_master_readdatavalid                       : std_logic;                     -- mm_interconnect_0:vide_dma_controller_CITANJE_0_avalon_dma_master_readdatavalid -> vide_dma_controller_CITANJE_0:master_readdatavalid
	signal vide_dma_controller_citanje_0_avalon_dma_master_lock                                : std_logic;                     -- vide_dma_controller_CITANJE_0:master_arbiterlock -> mm_interconnect_0:vide_dma_controller_CITANJE_0_avalon_dma_master_lock
	signal dma_controller_upis_avalon_dma_master_waitrequest                                   : std_logic;                     -- mm_interconnect_0:DMA_CONTROLLER_UPIS_avalon_dma_master_waitrequest -> DMA_CONTROLLER_UPIS:master_waitrequest
	signal dma_controller_upis_avalon_dma_master_address                                       : std_logic_vector(31 downto 0); -- DMA_CONTROLLER_UPIS:master_address -> mm_interconnect_0:DMA_CONTROLLER_UPIS_avalon_dma_master_address
	signal dma_controller_upis_avalon_dma_master_write                                         : std_logic;                     -- DMA_CONTROLLER_UPIS:master_write -> mm_interconnect_0:DMA_CONTROLLER_UPIS_avalon_dma_master_write
	signal dma_controller_upis_avalon_dma_master_writedata                                     : std_logic_vector(15 downto 0); -- DMA_CONTROLLER_UPIS:master_writedata -> mm_interconnect_0:DMA_CONTROLLER_UPIS_avalon_dma_master_writedata
	signal hps_h2f_axi_master_awburst                                                          : std_logic_vector(1 downto 0);  -- hps:h2f_AWBURST -> mm_interconnect_0:hps_h2f_axi_master_awburst
	signal hps_h2f_axi_master_arlen                                                            : std_logic_vector(3 downto 0);  -- hps:h2f_ARLEN -> mm_interconnect_0:hps_h2f_axi_master_arlen
	signal hps_h2f_axi_master_wstrb                                                            : std_logic_vector(7 downto 0);  -- hps:h2f_WSTRB -> mm_interconnect_0:hps_h2f_axi_master_wstrb
	signal hps_h2f_axi_master_wready                                                           : std_logic;                     -- mm_interconnect_0:hps_h2f_axi_master_wready -> hps:h2f_WREADY
	signal hps_h2f_axi_master_rid                                                              : std_logic_vector(11 downto 0); -- mm_interconnect_0:hps_h2f_axi_master_rid -> hps:h2f_RID
	signal hps_h2f_axi_master_rready                                                           : std_logic;                     -- hps:h2f_RREADY -> mm_interconnect_0:hps_h2f_axi_master_rready
	signal hps_h2f_axi_master_awlen                                                            : std_logic_vector(3 downto 0);  -- hps:h2f_AWLEN -> mm_interconnect_0:hps_h2f_axi_master_awlen
	signal hps_h2f_axi_master_wid                                                              : std_logic_vector(11 downto 0); -- hps:h2f_WID -> mm_interconnect_0:hps_h2f_axi_master_wid
	signal hps_h2f_axi_master_arcache                                                          : std_logic_vector(3 downto 0);  -- hps:h2f_ARCACHE -> mm_interconnect_0:hps_h2f_axi_master_arcache
	signal hps_h2f_axi_master_wvalid                                                           : std_logic;                     -- hps:h2f_WVALID -> mm_interconnect_0:hps_h2f_axi_master_wvalid
	signal hps_h2f_axi_master_araddr                                                           : std_logic_vector(29 downto 0); -- hps:h2f_ARADDR -> mm_interconnect_0:hps_h2f_axi_master_araddr
	signal hps_h2f_axi_master_arprot                                                           : std_logic_vector(2 downto 0);  -- hps:h2f_ARPROT -> mm_interconnect_0:hps_h2f_axi_master_arprot
	signal hps_h2f_axi_master_awprot                                                           : std_logic_vector(2 downto 0);  -- hps:h2f_AWPROT -> mm_interconnect_0:hps_h2f_axi_master_awprot
	signal hps_h2f_axi_master_wdata                                                            : std_logic_vector(63 downto 0); -- hps:h2f_WDATA -> mm_interconnect_0:hps_h2f_axi_master_wdata
	signal hps_h2f_axi_master_arvalid                                                          : std_logic;                     -- hps:h2f_ARVALID -> mm_interconnect_0:hps_h2f_axi_master_arvalid
	signal hps_h2f_axi_master_awcache                                                          : std_logic_vector(3 downto 0);  -- hps:h2f_AWCACHE -> mm_interconnect_0:hps_h2f_axi_master_awcache
	signal hps_h2f_axi_master_arid                                                             : std_logic_vector(11 downto 0); -- hps:h2f_ARID -> mm_interconnect_0:hps_h2f_axi_master_arid
	signal hps_h2f_axi_master_arlock                                                           : std_logic_vector(1 downto 0);  -- hps:h2f_ARLOCK -> mm_interconnect_0:hps_h2f_axi_master_arlock
	signal hps_h2f_axi_master_awlock                                                           : std_logic_vector(1 downto 0);  -- hps:h2f_AWLOCK -> mm_interconnect_0:hps_h2f_axi_master_awlock
	signal hps_h2f_axi_master_awaddr                                                           : std_logic_vector(29 downto 0); -- hps:h2f_AWADDR -> mm_interconnect_0:hps_h2f_axi_master_awaddr
	signal hps_h2f_axi_master_bresp                                                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hps_h2f_axi_master_bresp -> hps:h2f_BRESP
	signal hps_h2f_axi_master_arready                                                          : std_logic;                     -- mm_interconnect_0:hps_h2f_axi_master_arready -> hps:h2f_ARREADY
	signal hps_h2f_axi_master_rdata                                                            : std_logic_vector(63 downto 0); -- mm_interconnect_0:hps_h2f_axi_master_rdata -> hps:h2f_RDATA
	signal hps_h2f_axi_master_awready                                                          : std_logic;                     -- mm_interconnect_0:hps_h2f_axi_master_awready -> hps:h2f_AWREADY
	signal hps_h2f_axi_master_arburst                                                          : std_logic_vector(1 downto 0);  -- hps:h2f_ARBURST -> mm_interconnect_0:hps_h2f_axi_master_arburst
	signal hps_h2f_axi_master_arsize                                                           : std_logic_vector(2 downto 0);  -- hps:h2f_ARSIZE -> mm_interconnect_0:hps_h2f_axi_master_arsize
	signal hps_h2f_axi_master_bready                                                           : std_logic;                     -- hps:h2f_BREADY -> mm_interconnect_0:hps_h2f_axi_master_bready
	signal hps_h2f_axi_master_rlast                                                            : std_logic;                     -- mm_interconnect_0:hps_h2f_axi_master_rlast -> hps:h2f_RLAST
	signal hps_h2f_axi_master_wlast                                                            : std_logic;                     -- hps:h2f_WLAST -> mm_interconnect_0:hps_h2f_axi_master_wlast
	signal hps_h2f_axi_master_rresp                                                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hps_h2f_axi_master_rresp -> hps:h2f_RRESP
	signal hps_h2f_axi_master_awid                                                             : std_logic_vector(11 downto 0); -- hps:h2f_AWID -> mm_interconnect_0:hps_h2f_axi_master_awid
	signal hps_h2f_axi_master_bid                                                              : std_logic_vector(11 downto 0); -- mm_interconnect_0:hps_h2f_axi_master_bid -> hps:h2f_BID
	signal hps_h2f_axi_master_bvalid                                                           : std_logic;                     -- mm_interconnect_0:hps_h2f_axi_master_bvalid -> hps:h2f_BVALID
	signal hps_h2f_axi_master_awsize                                                           : std_logic_vector(2 downto 0);  -- hps:h2f_AWSIZE -> mm_interconnect_0:hps_h2f_axi_master_awsize
	signal hps_h2f_axi_master_awvalid                                                          : std_logic;                     -- hps:h2f_AWVALID -> mm_interconnect_0:hps_h2f_axi_master_awvalid
	signal hps_h2f_axi_master_rvalid                                                           : std_logic;                     -- mm_interconnect_0:hps_h2f_axi_master_rvalid -> hps:h2f_RVALID
	signal dma_afina_matrica_citanje_avalon_dma_master_waitrequest                             : std_logic;                     -- mm_interconnect_0:dma_afina_matrica_citanje_avalon_dma_master_waitrequest -> dma_afina_matrica_citanje:master_waitrequest
	signal dma_afina_matrica_citanje_avalon_dma_master_readdata                                : std_logic_vector(63 downto 0); -- mm_interconnect_0:dma_afina_matrica_citanje_avalon_dma_master_readdata -> dma_afina_matrica_citanje:master_readdata
	signal dma_afina_matrica_citanje_avalon_dma_master_address                                 : std_logic_vector(31 downto 0); -- dma_afina_matrica_citanje:master_address -> mm_interconnect_0:dma_afina_matrica_citanje_avalon_dma_master_address
	signal dma_afina_matrica_citanje_avalon_dma_master_read                                    : std_logic;                     -- dma_afina_matrica_citanje:master_read -> mm_interconnect_0:dma_afina_matrica_citanje_avalon_dma_master_read
	signal dma_afina_matrica_citanje_avalon_dma_master_readdatavalid                           : std_logic;                     -- mm_interconnect_0:dma_afina_matrica_citanje_avalon_dma_master_readdatavalid -> dma_afina_matrica_citanje:master_readdatavalid
	signal dma_afina_matrica_citanje_avalon_dma_master_lock                                    : std_logic;                     -- dma_afina_matrica_citanje:master_arbiterlock -> mm_interconnect_0:dma_afina_matrica_citanje_avalon_dma_master_lock
	signal mm_interconnect_0_sdram_controller_s1_chipselect                                    : std_logic;                     -- mm_interconnect_0:sdram_controller_s1_chipselect -> sdram_controller:az_cs
	signal mm_interconnect_0_sdram_controller_s1_readdata                                      : std_logic_vector(15 downto 0); -- sdram_controller:za_data -> mm_interconnect_0:sdram_controller_s1_readdata
	signal mm_interconnect_0_sdram_controller_s1_waitrequest                                   : std_logic;                     -- sdram_controller:za_waitrequest -> mm_interconnect_0:sdram_controller_s1_waitrequest
	signal mm_interconnect_0_sdram_controller_s1_address                                       : std_logic_vector(24 downto 0); -- mm_interconnect_0:sdram_controller_s1_address -> sdram_controller:az_addr
	signal mm_interconnect_0_sdram_controller_s1_read                                          : std_logic;                     -- mm_interconnect_0:sdram_controller_s1_read -> mm_interconnect_0_sdram_controller_s1_read:in
	signal mm_interconnect_0_sdram_controller_s1_byteenable                                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_controller_s1_byteenable -> mm_interconnect_0_sdram_controller_s1_byteenable:in
	signal mm_interconnect_0_sdram_controller_s1_readdatavalid                                 : std_logic;                     -- sdram_controller:za_valid -> mm_interconnect_0:sdram_controller_s1_readdatavalid
	signal mm_interconnect_0_sdram_controller_s1_write                                         : std_logic;                     -- mm_interconnect_0:sdram_controller_s1_write -> mm_interconnect_0_sdram_controller_s1_write:in
	signal mm_interconnect_0_sdram_controller_s1_writedata                                     : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_controller_s1_writedata -> sdram_controller:az_data
	signal mm_interconnect_0_affine_matrix_s1_chipselect                                       : std_logic;                     -- mm_interconnect_0:affine_matrix_s1_chipselect -> affine_matrix:chipselect
	signal mm_interconnect_0_affine_matrix_s1_readdata                                         : std_logic_vector(31 downto 0); -- affine_matrix:readdata -> mm_interconnect_0:affine_matrix_s1_readdata
	signal mm_interconnect_0_affine_matrix_s1_address                                          : std_logic_vector(9 downto 0);  -- mm_interconnect_0:affine_matrix_s1_address -> affine_matrix:address
	signal mm_interconnect_0_affine_matrix_s1_byteenable                                       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:affine_matrix_s1_byteenable -> affine_matrix:byteenable
	signal mm_interconnect_0_affine_matrix_s1_write                                            : std_logic;                     -- mm_interconnect_0:affine_matrix_s1_write -> affine_matrix:write
	signal mm_interconnect_0_affine_matrix_s1_writedata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:affine_matrix_s1_writedata -> affine_matrix:writedata
	signal mm_interconnect_0_affine_matrix_s1_clken                                            : std_logic;                     -- mm_interconnect_0:affine_matrix_s1_clken -> affine_matrix:clken
	signal hps_h2f_lw_axi_master_awburst                                                       : std_logic_vector(1 downto 0);  -- hps:h2f_lw_AWBURST -> mm_interconnect_1:hps_h2f_lw_axi_master_awburst
	signal hps_h2f_lw_axi_master_arlen                                                         : std_logic_vector(3 downto 0);  -- hps:h2f_lw_ARLEN -> mm_interconnect_1:hps_h2f_lw_axi_master_arlen
	signal hps_h2f_lw_axi_master_wstrb                                                         : std_logic_vector(3 downto 0);  -- hps:h2f_lw_WSTRB -> mm_interconnect_1:hps_h2f_lw_axi_master_wstrb
	signal hps_h2f_lw_axi_master_wready                                                        : std_logic;                     -- mm_interconnect_1:hps_h2f_lw_axi_master_wready -> hps:h2f_lw_WREADY
	signal hps_h2f_lw_axi_master_rid                                                           : std_logic_vector(11 downto 0); -- mm_interconnect_1:hps_h2f_lw_axi_master_rid -> hps:h2f_lw_RID
	signal hps_h2f_lw_axi_master_rready                                                        : std_logic;                     -- hps:h2f_lw_RREADY -> mm_interconnect_1:hps_h2f_lw_axi_master_rready
	signal hps_h2f_lw_axi_master_awlen                                                         : std_logic_vector(3 downto 0);  -- hps:h2f_lw_AWLEN -> mm_interconnect_1:hps_h2f_lw_axi_master_awlen
	signal hps_h2f_lw_axi_master_wid                                                           : std_logic_vector(11 downto 0); -- hps:h2f_lw_WID -> mm_interconnect_1:hps_h2f_lw_axi_master_wid
	signal hps_h2f_lw_axi_master_arcache                                                       : std_logic_vector(3 downto 0);  -- hps:h2f_lw_ARCACHE -> mm_interconnect_1:hps_h2f_lw_axi_master_arcache
	signal hps_h2f_lw_axi_master_wvalid                                                        : std_logic;                     -- hps:h2f_lw_WVALID -> mm_interconnect_1:hps_h2f_lw_axi_master_wvalid
	signal hps_h2f_lw_axi_master_araddr                                                        : std_logic_vector(20 downto 0); -- hps:h2f_lw_ARADDR -> mm_interconnect_1:hps_h2f_lw_axi_master_araddr
	signal hps_h2f_lw_axi_master_arprot                                                        : std_logic_vector(2 downto 0);  -- hps:h2f_lw_ARPROT -> mm_interconnect_1:hps_h2f_lw_axi_master_arprot
	signal hps_h2f_lw_axi_master_awprot                                                        : std_logic_vector(2 downto 0);  -- hps:h2f_lw_AWPROT -> mm_interconnect_1:hps_h2f_lw_axi_master_awprot
	signal hps_h2f_lw_axi_master_wdata                                                         : std_logic_vector(31 downto 0); -- hps:h2f_lw_WDATA -> mm_interconnect_1:hps_h2f_lw_axi_master_wdata
	signal hps_h2f_lw_axi_master_arvalid                                                       : std_logic;                     -- hps:h2f_lw_ARVALID -> mm_interconnect_1:hps_h2f_lw_axi_master_arvalid
	signal hps_h2f_lw_axi_master_awcache                                                       : std_logic_vector(3 downto 0);  -- hps:h2f_lw_AWCACHE -> mm_interconnect_1:hps_h2f_lw_axi_master_awcache
	signal hps_h2f_lw_axi_master_arid                                                          : std_logic_vector(11 downto 0); -- hps:h2f_lw_ARID -> mm_interconnect_1:hps_h2f_lw_axi_master_arid
	signal hps_h2f_lw_axi_master_arlock                                                        : std_logic_vector(1 downto 0);  -- hps:h2f_lw_ARLOCK -> mm_interconnect_1:hps_h2f_lw_axi_master_arlock
	signal hps_h2f_lw_axi_master_awlock                                                        : std_logic_vector(1 downto 0);  -- hps:h2f_lw_AWLOCK -> mm_interconnect_1:hps_h2f_lw_axi_master_awlock
	signal hps_h2f_lw_axi_master_awaddr                                                        : std_logic_vector(20 downto 0); -- hps:h2f_lw_AWADDR -> mm_interconnect_1:hps_h2f_lw_axi_master_awaddr
	signal hps_h2f_lw_axi_master_bresp                                                         : std_logic_vector(1 downto 0);  -- mm_interconnect_1:hps_h2f_lw_axi_master_bresp -> hps:h2f_lw_BRESP
	signal hps_h2f_lw_axi_master_arready                                                       : std_logic;                     -- mm_interconnect_1:hps_h2f_lw_axi_master_arready -> hps:h2f_lw_ARREADY
	signal hps_h2f_lw_axi_master_rdata                                                         : std_logic_vector(31 downto 0); -- mm_interconnect_1:hps_h2f_lw_axi_master_rdata -> hps:h2f_lw_RDATA
	signal hps_h2f_lw_axi_master_awready                                                       : std_logic;                     -- mm_interconnect_1:hps_h2f_lw_axi_master_awready -> hps:h2f_lw_AWREADY
	signal hps_h2f_lw_axi_master_arburst                                                       : std_logic_vector(1 downto 0);  -- hps:h2f_lw_ARBURST -> mm_interconnect_1:hps_h2f_lw_axi_master_arburst
	signal hps_h2f_lw_axi_master_arsize                                                        : std_logic_vector(2 downto 0);  -- hps:h2f_lw_ARSIZE -> mm_interconnect_1:hps_h2f_lw_axi_master_arsize
	signal hps_h2f_lw_axi_master_bready                                                        : std_logic;                     -- hps:h2f_lw_BREADY -> mm_interconnect_1:hps_h2f_lw_axi_master_bready
	signal hps_h2f_lw_axi_master_rlast                                                         : std_logic;                     -- mm_interconnect_1:hps_h2f_lw_axi_master_rlast -> hps:h2f_lw_RLAST
	signal hps_h2f_lw_axi_master_wlast                                                         : std_logic;                     -- hps:h2f_lw_WLAST -> mm_interconnect_1:hps_h2f_lw_axi_master_wlast
	signal hps_h2f_lw_axi_master_rresp                                                         : std_logic_vector(1 downto 0);  -- mm_interconnect_1:hps_h2f_lw_axi_master_rresp -> hps:h2f_lw_RRESP
	signal hps_h2f_lw_axi_master_awid                                                          : std_logic_vector(11 downto 0); -- hps:h2f_lw_AWID -> mm_interconnect_1:hps_h2f_lw_axi_master_awid
	signal hps_h2f_lw_axi_master_bid                                                           : std_logic_vector(11 downto 0); -- mm_interconnect_1:hps_h2f_lw_axi_master_bid -> hps:h2f_lw_BID
	signal hps_h2f_lw_axi_master_bvalid                                                        : std_logic;                     -- mm_interconnect_1:hps_h2f_lw_axi_master_bvalid -> hps:h2f_lw_BVALID
	signal hps_h2f_lw_axi_master_awsize                                                        : std_logic_vector(2 downto 0);  -- hps:h2f_lw_AWSIZE -> mm_interconnect_1:hps_h2f_lw_axi_master_awsize
	signal hps_h2f_lw_axi_master_awvalid                                                       : std_logic;                     -- hps:h2f_lw_AWVALID -> mm_interconnect_1:hps_h2f_lw_axi_master_awvalid
	signal hps_h2f_lw_axi_master_rvalid                                                        : std_logic;                     -- mm_interconnect_1:hps_h2f_lw_axi_master_rvalid -> hps:h2f_lw_RVALID
	signal mm_interconnect_1_vide_dma_controller_avalon_dma_control_slave_readdata             : std_logic_vector(31 downto 0); -- vide_dma_controller:slave_readdata -> mm_interconnect_1:vide_dma_controller_avalon_dma_control_slave_readdata
	signal mm_interconnect_1_vide_dma_controller_avalon_dma_control_slave_address              : std_logic_vector(1 downto 0);  -- mm_interconnect_1:vide_dma_controller_avalon_dma_control_slave_address -> vide_dma_controller:slave_address
	signal mm_interconnect_1_vide_dma_controller_avalon_dma_control_slave_read                 : std_logic;                     -- mm_interconnect_1:vide_dma_controller_avalon_dma_control_slave_read -> vide_dma_controller:slave_read
	signal mm_interconnect_1_vide_dma_controller_avalon_dma_control_slave_byteenable           : std_logic_vector(3 downto 0);  -- mm_interconnect_1:vide_dma_controller_avalon_dma_control_slave_byteenable -> vide_dma_controller:slave_byteenable
	signal mm_interconnect_1_vide_dma_controller_avalon_dma_control_slave_write                : std_logic;                     -- mm_interconnect_1:vide_dma_controller_avalon_dma_control_slave_write -> vide_dma_controller:slave_write
	signal mm_interconnect_1_vide_dma_controller_avalon_dma_control_slave_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_1:vide_dma_controller_avalon_dma_control_slave_writedata -> vide_dma_controller:slave_writedata
	signal mm_interconnect_1_vide_dma_controller_citanje_avalon_dma_control_slave_readdata     : std_logic_vector(31 downto 0); -- vide_dma_controller_CITANJE:slave_readdata -> mm_interconnect_1:vide_dma_controller_CITANJE_avalon_dma_control_slave_readdata
	signal mm_interconnect_1_vide_dma_controller_citanje_avalon_dma_control_slave_address      : std_logic_vector(1 downto 0);  -- mm_interconnect_1:vide_dma_controller_CITANJE_avalon_dma_control_slave_address -> vide_dma_controller_CITANJE:slave_address
	signal mm_interconnect_1_vide_dma_controller_citanje_avalon_dma_control_slave_read         : std_logic;                     -- mm_interconnect_1:vide_dma_controller_CITANJE_avalon_dma_control_slave_read -> vide_dma_controller_CITANJE:slave_read
	signal mm_interconnect_1_vide_dma_controller_citanje_avalon_dma_control_slave_byteenable   : std_logic_vector(3 downto 0);  -- mm_interconnect_1:vide_dma_controller_CITANJE_avalon_dma_control_slave_byteenable -> vide_dma_controller_CITANJE:slave_byteenable
	signal mm_interconnect_1_vide_dma_controller_citanje_avalon_dma_control_slave_write        : std_logic;                     -- mm_interconnect_1:vide_dma_controller_CITANJE_avalon_dma_control_slave_write -> vide_dma_controller_CITANJE:slave_write
	signal mm_interconnect_1_vide_dma_controller_citanje_avalon_dma_control_slave_writedata    : std_logic_vector(31 downto 0); -- mm_interconnect_1:vide_dma_controller_CITANJE_avalon_dma_control_slave_writedata -> vide_dma_controller_CITANJE:slave_writedata
	signal mm_interconnect_1_dma_controller_upis_avalon_dma_control_slave_readdata             : std_logic_vector(31 downto 0); -- DMA_CONTROLLER_UPIS:slave_readdata -> mm_interconnect_1:DMA_CONTROLLER_UPIS_avalon_dma_control_slave_readdata
	signal mm_interconnect_1_dma_controller_upis_avalon_dma_control_slave_address              : std_logic_vector(1 downto 0);  -- mm_interconnect_1:DMA_CONTROLLER_UPIS_avalon_dma_control_slave_address -> DMA_CONTROLLER_UPIS:slave_address
	signal mm_interconnect_1_dma_controller_upis_avalon_dma_control_slave_read                 : std_logic;                     -- mm_interconnect_1:DMA_CONTROLLER_UPIS_avalon_dma_control_slave_read -> DMA_CONTROLLER_UPIS:slave_read
	signal mm_interconnect_1_dma_controller_upis_avalon_dma_control_slave_byteenable           : std_logic_vector(3 downto 0);  -- mm_interconnect_1:DMA_CONTROLLER_UPIS_avalon_dma_control_slave_byteenable -> DMA_CONTROLLER_UPIS:slave_byteenable
	signal mm_interconnect_1_dma_controller_upis_avalon_dma_control_slave_write                : std_logic;                     -- mm_interconnect_1:DMA_CONTROLLER_UPIS_avalon_dma_control_slave_write -> DMA_CONTROLLER_UPIS:slave_write
	signal mm_interconnect_1_dma_controller_upis_avalon_dma_control_slave_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_1:DMA_CONTROLLER_UPIS_avalon_dma_control_slave_writedata -> DMA_CONTROLLER_UPIS:slave_writedata
	signal mm_interconnect_1_vide_dma_controller_citanje_0_avalon_dma_control_slave_readdata   : std_logic_vector(31 downto 0); -- vide_dma_controller_CITANJE_0:slave_readdata -> mm_interconnect_1:vide_dma_controller_CITANJE_0_avalon_dma_control_slave_readdata
	signal mm_interconnect_1_vide_dma_controller_citanje_0_avalon_dma_control_slave_address    : std_logic_vector(1 downto 0);  -- mm_interconnect_1:vide_dma_controller_CITANJE_0_avalon_dma_control_slave_address -> vide_dma_controller_CITANJE_0:slave_address
	signal mm_interconnect_1_vide_dma_controller_citanje_0_avalon_dma_control_slave_read       : std_logic;                     -- mm_interconnect_1:vide_dma_controller_CITANJE_0_avalon_dma_control_slave_read -> vide_dma_controller_CITANJE_0:slave_read
	signal mm_interconnect_1_vide_dma_controller_citanje_0_avalon_dma_control_slave_byteenable : std_logic_vector(3 downto 0);  -- mm_interconnect_1:vide_dma_controller_CITANJE_0_avalon_dma_control_slave_byteenable -> vide_dma_controller_CITANJE_0:slave_byteenable
	signal mm_interconnect_1_vide_dma_controller_citanje_0_avalon_dma_control_slave_write      : std_logic;                     -- mm_interconnect_1:vide_dma_controller_CITANJE_0_avalon_dma_control_slave_write -> vide_dma_controller_CITANJE_0:slave_write
	signal mm_interconnect_1_vide_dma_controller_citanje_0_avalon_dma_control_slave_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_1:vide_dma_controller_CITANJE_0_avalon_dma_control_slave_writedata -> vide_dma_controller_CITANJE_0:slave_writedata
	signal mm_interconnect_1_izbor_prikaza_slike_0_izbor_slike_readdata                        : std_logic_vector(31 downto 0); -- Izbor_Prikaza_Slike_0:izbor_slike_readdata -> mm_interconnect_1:Izbor_Prikaza_Slike_0_izbor_slike_readdata
	signal mm_interconnect_1_izbor_prikaza_slike_0_izbor_slike_address                         : std_logic_vector(7 downto 0);  -- mm_interconnect_1:Izbor_Prikaza_Slike_0_izbor_slike_address -> Izbor_Prikaza_Slike_0:izbor_slike_address
	signal mm_interconnect_1_izbor_prikaza_slike_0_izbor_slike_read                            : std_logic;                     -- mm_interconnect_1:Izbor_Prikaza_Slike_0_izbor_slike_read -> Izbor_Prikaza_Slike_0:izbor_slike_read
	signal mm_interconnect_1_izbor_prikaza_slike_0_izbor_slike_write                           : std_logic;                     -- mm_interconnect_1:Izbor_Prikaza_Slike_0_izbor_slike_write -> Izbor_Prikaza_Slike_0:izbor_slike_write
	signal mm_interconnect_1_izbor_prikaza_slike_0_izbor_slike_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_1:Izbor_Prikaza_Slike_0_izbor_slike_writedata -> Izbor_Prikaza_Slike_0:izbor_slike_writedata
	signal mm_interconnect_1_image_processing_0_s0_readdata                                    : std_logic_vector(31 downto 0); -- Image_Processing_0:avs_s0_readdata -> mm_interconnect_1:Image_Processing_0_s0_readdata
	signal mm_interconnect_1_image_processing_0_s0_address                                     : std_logic_vector(7 downto 0);  -- mm_interconnect_1:Image_Processing_0_s0_address -> Image_Processing_0:avs_s0_address
	signal mm_interconnect_1_image_processing_0_s0_read                                        : std_logic;                     -- mm_interconnect_1:Image_Processing_0_s0_read -> Image_Processing_0:avs_s0_read
	signal mm_interconnect_1_image_processing_0_s0_write                                       : std_logic;                     -- mm_interconnect_1:Image_Processing_0_s0_write -> Image_Processing_0:avs_s0_write
	signal mm_interconnect_1_image_processing_0_s0_writedata                                   : std_logic_vector(31 downto 0); -- mm_interconnect_1:Image_Processing_0_s0_writedata -> Image_Processing_0:avs_s0_writedata
	signal izbor_prikaza_slike_0_led_master_waitrequest                                        : std_logic;                     -- mm_interconnect_2:Izbor_Prikaza_Slike_0_led_master_waitrequest -> Izbor_Prikaza_Slike_0:led_master_waitrequest
	signal izbor_prikaza_slike_0_led_master_write                                              : std_logic;                     -- Izbor_Prikaza_Slike_0:led_master_write -> mm_interconnect_2:Izbor_Prikaza_Slike_0_led_master_write
	signal izbor_prikaza_slike_0_led_master_writedata                                          : std_logic_vector(7 downto 0);  -- Izbor_Prikaza_Slike_0:led_master_writedata -> mm_interconnect_2:Izbor_Prikaza_Slike_0_led_master_writedata
	signal mm_interconnect_2_led_indication_0_s1_chipselect                                    : std_logic;                     -- mm_interconnect_2:led_indication_0_s1_chipselect -> led_indication_0:chipselect
	signal mm_interconnect_2_led_indication_0_s1_readdata                                      : std_logic_vector(31 downto 0); -- led_indication_0:readdata -> mm_interconnect_2:led_indication_0_s1_readdata
	signal mm_interconnect_2_led_indication_0_s1_address                                       : std_logic_vector(1 downto 0);  -- mm_interconnect_2:led_indication_0_s1_address -> led_indication_0:address
	signal mm_interconnect_2_led_indication_0_s1_write                                         : std_logic;                     -- mm_interconnect_2:led_indication_0_s1_write -> mm_interconnect_2_led_indication_0_s1_write:in
	signal mm_interconnect_2_led_indication_0_s1_writedata                                     : std_logic_vector(31 downto 0); -- mm_interconnect_2:led_indication_0_s1_writedata -> led_indication_0:writedata
	signal rst_controller_reset_out_reset                                                      : std_logic;                     -- rst_controller:reset_out -> [DMA_CONTROLLER_UPIS:reset, Image_Processing_0:reset_reset, Izbor_Prikaza_Slike_0:reset_reset, Pozicioniranje_Piksela_u_SDRAM_0:reset_reset, Transformacija_Pozicije_Piksela:reset_reset, affine_matrix:reset, affine_matrix:reset2, dma_afina_matrica_citanje:reset, mm_interconnect_0:vide_dma_controller_reset_reset_bridge_in_reset_reset, mm_interconnect_1:vide_dma_controller_reset_reset_bridge_in_reset_reset, mm_interconnect_2:Izbor_Prikaza_Slike_0_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset, vide_dma_controller:reset, vide_dma_controller_CITANJE:reset, vide_dma_controller_CITANJE_0:reset, video_dual_clock_buffer:reset_stream_in]
	signal rst_controller_reset_out_reset_req                                                  : std_logic;                     -- rst_controller:reset_req -> [affine_matrix:reset_req, affine_matrix:reset_req2, rst_translator:reset_req_in]
	signal rst_controller_001_reset_out_reset                                                  : std_logic;                     -- rst_controller_001:reset_out -> [video_dual_clock_buffer:reset_stream_out, video_rgb_resampler_0:reset, video_vga_controller:reset]
	signal rst_controller_002_reset_out_reset                                                  : std_logic;                     -- rst_controller_002:reset_out -> [mm_interconnect_0:hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]
	signal hps_h2f_reset_reset_ports_inv                                                       : std_logic;                     -- hps_h2f_reset_reset:inv -> [rst_controller_002:reset_in0, sys_sdram_pll:ref_reset_reset]
	signal mm_interconnect_0_sdram_controller_s1_read_ports_inv                                : std_logic;                     -- mm_interconnect_0_sdram_controller_s1_read:inv -> sdram_controller:az_rd_n
	signal mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_controller_s1_byteenable:inv -> sdram_controller:az_be_n
	signal mm_interconnect_0_sdram_controller_s1_write_ports_inv                               : std_logic;                     -- mm_interconnect_0_sdram_controller_s1_write:inv -> sdram_controller:az_wr_n
	signal mm_interconnect_2_led_indication_0_s1_write_ports_inv                               : std_logic;                     -- mm_interconnect_2_led_indication_0_s1_write:inv -> led_indication_0:write_n
	signal rst_controller_reset_out_reset_ports_inv                                            : std_logic;                     -- rst_controller_reset_out_reset:inv -> [led_indication_0:reset_n, sdram_controller:reset_n]

begin

	dma_controller_upis : component VideoBox_DMA_CONTROLLER_UPIS
		port map (
			clk                  => sys_sdram_pll_sys_clk_clk,                                                 --                      clk.clk
			reset                => rst_controller_reset_out_reset,                                            --                    reset.reset
			stream_data          => image_processing_0_out0_data,                                              --          avalon_dma_sink.data
			stream_startofpacket => image_processing_0_out0_startofpacket,                                     --                         .startofpacket
			stream_endofpacket   => image_processing_0_out0_endofpacket,                                       --                         .endofpacket
			stream_valid         => image_processing_0_out0_valid,                                             --                         .valid
			stream_ready         => image_processing_0_out0_ready,                                             --                         .ready
			slave_address        => mm_interconnect_1_dma_controller_upis_avalon_dma_control_slave_address,    -- avalon_dma_control_slave.address
			slave_byteenable     => mm_interconnect_1_dma_controller_upis_avalon_dma_control_slave_byteenable, --                         .byteenable
			slave_read           => mm_interconnect_1_dma_controller_upis_avalon_dma_control_slave_read,       --                         .read
			slave_write          => mm_interconnect_1_dma_controller_upis_avalon_dma_control_slave_write,      --                         .write
			slave_writedata      => mm_interconnect_1_dma_controller_upis_avalon_dma_control_slave_writedata,  --                         .writedata
			slave_readdata       => mm_interconnect_1_dma_controller_upis_avalon_dma_control_slave_readdata,   --                         .readdata
			master_address       => dma_controller_upis_avalon_dma_master_address,                             --        avalon_dma_master.address
			master_waitrequest   => dma_controller_upis_avalon_dma_master_waitrequest,                         --                         .waitrequest
			master_write         => dma_controller_upis_avalon_dma_master_write,                               --                         .write
			master_writedata     => dma_controller_upis_avalon_dma_master_writedata                            --                         .writedata
		);

	image_processing_0 : component Image_Processing
		port map (
			avs_s0_address         => mm_interconnect_1_image_processing_0_s0_address,                 --    s0.address
			avs_s0_read            => mm_interconnect_1_image_processing_0_s0_read,                    --      .read
			avs_s0_readdata        => mm_interconnect_1_image_processing_0_s0_readdata,                --      .readdata
			avs_s0_write           => mm_interconnect_1_image_processing_0_s0_write,                   --      .write
			avs_s0_writedata       => mm_interconnect_1_image_processing_0_s0_writedata,               --      .writedata
			asi_in0_data           => vide_dma_controller_citanje_0_avalon_pixel_source_data,          --   in0.data
			asi_in0_ready          => vide_dma_controller_citanje_0_avalon_pixel_source_ready,         --      .ready
			asi_in0_valid          => vide_dma_controller_citanje_0_avalon_pixel_source_valid,         --      .valid
			asi_in0_endofpacket    => vide_dma_controller_citanje_0_avalon_pixel_source_endofpacket,   --      .endofpacket
			asi_in0_startofpacket  => vide_dma_controller_citanje_0_avalon_pixel_source_startofpacket, --      .startofpacket
			aso_out0_data          => image_processing_0_out0_data,                                    --  out0.data
			aso_out0_ready         => image_processing_0_out0_ready,                                   --      .ready
			aso_out0_valid         => image_processing_0_out0_valid,                                   --      .valid
			aso_out0_endofpacket   => image_processing_0_out0_endofpacket,                             --      .endofpacket
			aso_out0_startofpacket => image_processing_0_out0_startofpacket,                           --      .startofpacket
			reset_reset            => rst_controller_reset_out_reset,                                  -- reset.reset
			clock_clk              => sys_sdram_pll_sys_clk_clk                                        -- clock.clk
		);

	izbor_prikaza_slike_0 : component Izbor_Prikaza_Slike
		port map (
			out_data               => izbor_prikaza_slike_0_out_data,                                --         out.data
			out_endofpacket        => izbor_prikaza_slike_0_out_endofpacket,                         --            .endofpacket
			out_ready              => izbor_prikaza_slike_0_out_ready,                               --            .ready
			out_startofpacket      => izbor_prikaza_slike_0_out_startofpacket,                       --            .startofpacket
			out_valid              => izbor_prikaza_slike_0_out_valid,                               --            .valid
			in1_valid              => vide_dma_controller_citanje_avalon_pixel_source_valid,         --         in1.valid
			in1_startofpacket      => vide_dma_controller_citanje_avalon_pixel_source_startofpacket, --            .startofpacket
			in1_ready              => vide_dma_controller_citanje_avalon_pixel_source_ready,         --            .ready
			in1_endofpacket        => vide_dma_controller_citanje_avalon_pixel_source_endofpacket,   --            .endofpacket
			in1_data               => vide_dma_controller_citanje_avalon_pixel_source_data,          --            .data
			in2_data               => vide_dma_controller_avalon_pixel_source_data,                  --         in2.data
			in2_ready              => vide_dma_controller_avalon_pixel_source_ready,                 --            .ready
			in2_valid              => vide_dma_controller_avalon_pixel_source_valid,                 --            .valid
			in2_startofpacket      => vide_dma_controller_avalon_pixel_source_startofpacket,         --            .startofpacket
			in2_endofpacket        => vide_dma_controller_avalon_pixel_source_endofpacket,           --            .endofpacket
			clock_clk              => sys_sdram_pll_sys_clk_clk,                                     --       clock.clk
			reset_reset            => rst_controller_reset_out_reset,                                --       reset.reset
			izbor_slike_address    => mm_interconnect_1_izbor_prikaza_slike_0_izbor_slike_address,   -- izbor_slike.address
			izbor_slike_write      => mm_interconnect_1_izbor_prikaza_slike_0_izbor_slike_write,     --            .write
			izbor_slike_writedata  => mm_interconnect_1_izbor_prikaza_slike_0_izbor_slike_writedata, --            .writedata
			izbor_slike_read       => mm_interconnect_1_izbor_prikaza_slike_0_izbor_slike_read,      --            .read
			izbor_slike_readdata   => mm_interconnect_1_izbor_prikaza_slike_0_izbor_slike_readdata,  --            .readdata
			led_master_write       => izbor_prikaza_slike_0_led_master_write,                        --  led_master.write
			led_master_writedata   => izbor_prikaza_slike_0_led_master_writedata,                    --            .writedata
			led_master_waitrequest => izbor_prikaza_slike_0_led_master_waitrequest                   --            .waitrequest
		);

	pozicioniranje_piksela_u_sdram_0 : component Pozicioniranje_Piksela_u_SDRAM
		port map (
			reset_reset              => rst_controller_reset_out_reset,                       --      reset.reset
			clock_clk                => sys_sdram_pll_sys_clk_clk,                            --      clock.clk
			out_piksel_data          => open,                                                 -- out_piksel.data
			out_piksel_endofpacket   => open,                                                 --           .endofpacket
			out_piksel_ready         => open,                                                 --           .ready
			out_piksel_startofpacket => open,                                                 --           .startofpacket
			out_piksel_valid         => open,                                                 --           .valid
			in_piksel_ready          => open,                                                 --  in_piksel.ready
			in_piksel_valid          => open,                                                 --           .valid
			in_piksel_endofpacket    => open,                                                 --           .endofpacket
			in_piksel_data           => open,                                                 --           .data
			in_piksel_startofpacket  => open,                                                 --           .startofpacket
			in_xy_valid              => transformacija_pozicije_piksela_xy_out_valid,         --    in_xy_1.valid
			in_xy_startofpacket      => transformacija_pozicije_piksela_xy_out_startofpacket, --           .startofpacket
			in_xy_endofpacket        => transformacija_pozicije_piksela_xy_out_endofpacket,   --           .endofpacket
			in_xy_ready              => transformacija_pozicije_piksela_xy_out_ready,         --           .ready
			in_xy_data               => transformacija_pozicije_piksela_xy_out_data           --           .data
		);

	transformacija_pozicije_piksela : component Transformacija_Slike
		port map (
			clock_clk              => sys_sdram_pll_sys_clk_clk,                                   --                  clock.clk
			reset_reset            => rst_controller_reset_out_reset,                              --                  reset.reset
			out_data               => transformacija_pozicije_piksela_xy_out_data,                 --                 xy_out.data
			out_ready              => transformacija_pozicije_piksela_xy_out_ready,                --                       .ready
			out_startofpacket      => transformacija_pozicije_piksela_xy_out_startofpacket,        --                       .startofpacket
			out_endofpacket        => transformacija_pozicije_piksela_xy_out_endofpacket,          --                       .endofpacket
			out_valid              => transformacija_pozicije_piksela_xy_out_valid,                --                       .valid
			avalon_slave_write     => open,                                                        -- avalon_slave_parametar.write
			avalon_slave_writedata => open,                                                        --                       .writedata
			in_data                => dma_afina_matrica_citanje_avalon_pixel_source_data,          --          in_dma_affine.data
			in_ready               => dma_afina_matrica_citanje_avalon_pixel_source_ready,         --                       .ready
			in_startofpacket       => dma_afina_matrica_citanje_avalon_pixel_source_startofpacket, --                       .startofpacket
			in_endofpacket         => dma_afina_matrica_citanje_avalon_pixel_source_endofpacket,   --                       .endofpacket
			in_valid               => dma_afina_matrica_citanje_avalon_pixel_source_valid          --                       .valid
		);

	affine_matrix : component VideoBox_affine_matrix
		port map (
			clk         => sys_sdram_pll_sys_clk_clk,                     --   clk1.clk
			address     => mm_interconnect_0_affine_matrix_s1_address,    --     s1.address
			clken       => mm_interconnect_0_affine_matrix_s1_clken,      --       .clken
			chipselect  => mm_interconnect_0_affine_matrix_s1_chipselect, --       .chipselect
			write       => mm_interconnect_0_affine_matrix_s1_write,      --       .write
			readdata    => mm_interconnect_0_affine_matrix_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_0_affine_matrix_s1_writedata,  --       .writedata
			byteenable  => mm_interconnect_0_affine_matrix_s1_byteenable, --       .byteenable
			reset       => rst_controller_reset_out_reset,                -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,            --       .reset_req
			address2    => open,                                          --     s2.address
			chipselect2 => open,                                          --       .chipselect
			clken2      => open,                                          --       .clken
			write2      => open,                                          --       .write
			readdata2   => open,                                          --       .readdata
			writedata2  => open,                                          --       .writedata
			byteenable2 => open,                                          --       .byteenable
			clk2        => sys_sdram_pll_sys_clk_clk,                     --   clk2.clk
			reset2      => rst_controller_reset_out_reset,                -- reset2.reset
			reset_req2  => rst_controller_reset_out_reset_req,            --       .reset_req
			freeze      => '0'                                            -- (terminated)
		);

	dma_afina_matrica_citanje : component VideoBox_dma_afina_matrica_citanje
		port map (
			clk                  => sys_sdram_pll_sys_clk_clk,                                   --                      clk.clk
			reset                => rst_controller_reset_out_reset,                              --                    reset.reset
			master_address       => dma_afina_matrica_citanje_avalon_dma_master_address,         --        avalon_dma_master.address
			master_waitrequest   => dma_afina_matrica_citanje_avalon_dma_master_waitrequest,     --                         .waitrequest
			master_arbiterlock   => dma_afina_matrica_citanje_avalon_dma_master_lock,            --                         .lock
			master_read          => dma_afina_matrica_citanje_avalon_dma_master_read,            --                         .read
			master_readdata      => dma_afina_matrica_citanje_avalon_dma_master_readdata,        --                         .readdata
			master_readdatavalid => dma_afina_matrica_citanje_avalon_dma_master_readdatavalid,   --                         .readdatavalid
			slave_address        => open,                                                        -- avalon_dma_control_slave.address
			slave_byteenable     => open,                                                        --                         .byteenable
			slave_read           => open,                                                        --                         .read
			slave_write          => open,                                                        --                         .write
			slave_writedata      => open,                                                        --                         .writedata
			slave_readdata       => open,                                                        --                         .readdata
			stream_ready         => dma_afina_matrica_citanje_avalon_pixel_source_ready,         --      avalon_pixel_source.ready
			stream_data          => dma_afina_matrica_citanje_avalon_pixel_source_data,          --                         .data
			stream_startofpacket => dma_afina_matrica_citanje_avalon_pixel_source_startofpacket, --                         .startofpacket
			stream_endofpacket   => dma_afina_matrica_citanje_avalon_pixel_source_endofpacket,   --                         .endofpacket
			stream_valid         => dma_afina_matrica_citanje_avalon_pixel_source_valid          --                         .valid
		);

	hps : component VideoBox_hps
		generic map (
			F2S_Width => 0,
			S2F_Width => 2
		)
		port map (
			mem_a          => memory_mem_a,                  --            memory.mem_a
			mem_ba         => memory_mem_ba,                 --                  .mem_ba
			mem_ck         => memory_mem_ck,                 --                  .mem_ck
			mem_ck_n       => memory_mem_ck_n,               --                  .mem_ck_n
			mem_cke        => memory_mem_cke,                --                  .mem_cke
			mem_cs_n       => memory_mem_cs_n,               --                  .mem_cs_n
			mem_ras_n      => memory_mem_ras_n,              --                  .mem_ras_n
			mem_cas_n      => memory_mem_cas_n,              --                  .mem_cas_n
			mem_we_n       => memory_mem_we_n,               --                  .mem_we_n
			mem_reset_n    => memory_mem_reset_n,            --                  .mem_reset_n
			mem_dq         => memory_mem_dq,                 --                  .mem_dq
			mem_dqs        => memory_mem_dqs,                --                  .mem_dqs
			mem_dqs_n      => memory_mem_dqs_n,              --                  .mem_dqs_n
			mem_odt        => memory_mem_odt,                --                  .mem_odt
			mem_dm         => memory_mem_dm,                 --                  .mem_dm
			oct_rzqin      => memory_oct_rzqin,              --                  .oct_rzqin
			h2f_rst_n      => hps_h2f_reset_reset,           --         h2f_reset.reset_n
			h2f_axi_clk    => sys_sdram_pll_sys_clk_clk,     --     h2f_axi_clock.clk
			h2f_AWID       => hps_h2f_axi_master_awid,       --    h2f_axi_master.awid
			h2f_AWADDR     => hps_h2f_axi_master_awaddr,     --                  .awaddr
			h2f_AWLEN      => hps_h2f_axi_master_awlen,      --                  .awlen
			h2f_AWSIZE     => hps_h2f_axi_master_awsize,     --                  .awsize
			h2f_AWBURST    => hps_h2f_axi_master_awburst,    --                  .awburst
			h2f_AWLOCK     => hps_h2f_axi_master_awlock,     --                  .awlock
			h2f_AWCACHE    => hps_h2f_axi_master_awcache,    --                  .awcache
			h2f_AWPROT     => hps_h2f_axi_master_awprot,     --                  .awprot
			h2f_AWVALID    => hps_h2f_axi_master_awvalid,    --                  .awvalid
			h2f_AWREADY    => hps_h2f_axi_master_awready,    --                  .awready
			h2f_WID        => hps_h2f_axi_master_wid,        --                  .wid
			h2f_WDATA      => hps_h2f_axi_master_wdata,      --                  .wdata
			h2f_WSTRB      => hps_h2f_axi_master_wstrb,      --                  .wstrb
			h2f_WLAST      => hps_h2f_axi_master_wlast,      --                  .wlast
			h2f_WVALID     => hps_h2f_axi_master_wvalid,     --                  .wvalid
			h2f_WREADY     => hps_h2f_axi_master_wready,     --                  .wready
			h2f_BID        => hps_h2f_axi_master_bid,        --                  .bid
			h2f_BRESP      => hps_h2f_axi_master_bresp,      --                  .bresp
			h2f_BVALID     => hps_h2f_axi_master_bvalid,     --                  .bvalid
			h2f_BREADY     => hps_h2f_axi_master_bready,     --                  .bready
			h2f_ARID       => hps_h2f_axi_master_arid,       --                  .arid
			h2f_ARADDR     => hps_h2f_axi_master_araddr,     --                  .araddr
			h2f_ARLEN      => hps_h2f_axi_master_arlen,      --                  .arlen
			h2f_ARSIZE     => hps_h2f_axi_master_arsize,     --                  .arsize
			h2f_ARBURST    => hps_h2f_axi_master_arburst,    --                  .arburst
			h2f_ARLOCK     => hps_h2f_axi_master_arlock,     --                  .arlock
			h2f_ARCACHE    => hps_h2f_axi_master_arcache,    --                  .arcache
			h2f_ARPROT     => hps_h2f_axi_master_arprot,     --                  .arprot
			h2f_ARVALID    => hps_h2f_axi_master_arvalid,    --                  .arvalid
			h2f_ARREADY    => hps_h2f_axi_master_arready,    --                  .arready
			h2f_RID        => hps_h2f_axi_master_rid,        --                  .rid
			h2f_RDATA      => hps_h2f_axi_master_rdata,      --                  .rdata
			h2f_RRESP      => hps_h2f_axi_master_rresp,      --                  .rresp
			h2f_RLAST      => hps_h2f_axi_master_rlast,      --                  .rlast
			h2f_RVALID     => hps_h2f_axi_master_rvalid,     --                  .rvalid
			h2f_RREADY     => hps_h2f_axi_master_rready,     --                  .rready
			h2f_lw_axi_clk => sys_sdram_pll_sys_clk_clk,     --  h2f_lw_axi_clock.clk
			h2f_lw_AWID    => hps_h2f_lw_axi_master_awid,    -- h2f_lw_axi_master.awid
			h2f_lw_AWADDR  => hps_h2f_lw_axi_master_awaddr,  --                  .awaddr
			h2f_lw_AWLEN   => hps_h2f_lw_axi_master_awlen,   --                  .awlen
			h2f_lw_AWSIZE  => hps_h2f_lw_axi_master_awsize,  --                  .awsize
			h2f_lw_AWBURST => hps_h2f_lw_axi_master_awburst, --                  .awburst
			h2f_lw_AWLOCK  => hps_h2f_lw_axi_master_awlock,  --                  .awlock
			h2f_lw_AWCACHE => hps_h2f_lw_axi_master_awcache, --                  .awcache
			h2f_lw_AWPROT  => hps_h2f_lw_axi_master_awprot,  --                  .awprot
			h2f_lw_AWVALID => hps_h2f_lw_axi_master_awvalid, --                  .awvalid
			h2f_lw_AWREADY => hps_h2f_lw_axi_master_awready, --                  .awready
			h2f_lw_WID     => hps_h2f_lw_axi_master_wid,     --                  .wid
			h2f_lw_WDATA   => hps_h2f_lw_axi_master_wdata,   --                  .wdata
			h2f_lw_WSTRB   => hps_h2f_lw_axi_master_wstrb,   --                  .wstrb
			h2f_lw_WLAST   => hps_h2f_lw_axi_master_wlast,   --                  .wlast
			h2f_lw_WVALID  => hps_h2f_lw_axi_master_wvalid,  --                  .wvalid
			h2f_lw_WREADY  => hps_h2f_lw_axi_master_wready,  --                  .wready
			h2f_lw_BID     => hps_h2f_lw_axi_master_bid,     --                  .bid
			h2f_lw_BRESP   => hps_h2f_lw_axi_master_bresp,   --                  .bresp
			h2f_lw_BVALID  => hps_h2f_lw_axi_master_bvalid,  --                  .bvalid
			h2f_lw_BREADY  => hps_h2f_lw_axi_master_bready,  --                  .bready
			h2f_lw_ARID    => hps_h2f_lw_axi_master_arid,    --                  .arid
			h2f_lw_ARADDR  => hps_h2f_lw_axi_master_araddr,  --                  .araddr
			h2f_lw_ARLEN   => hps_h2f_lw_axi_master_arlen,   --                  .arlen
			h2f_lw_ARSIZE  => hps_h2f_lw_axi_master_arsize,  --                  .arsize
			h2f_lw_ARBURST => hps_h2f_lw_axi_master_arburst, --                  .arburst
			h2f_lw_ARLOCK  => hps_h2f_lw_axi_master_arlock,  --                  .arlock
			h2f_lw_ARCACHE => hps_h2f_lw_axi_master_arcache, --                  .arcache
			h2f_lw_ARPROT  => hps_h2f_lw_axi_master_arprot,  --                  .arprot
			h2f_lw_ARVALID => hps_h2f_lw_axi_master_arvalid, --                  .arvalid
			h2f_lw_ARREADY => hps_h2f_lw_axi_master_arready, --                  .arready
			h2f_lw_RID     => hps_h2f_lw_axi_master_rid,     --                  .rid
			h2f_lw_RDATA   => hps_h2f_lw_axi_master_rdata,   --                  .rdata
			h2f_lw_RRESP   => hps_h2f_lw_axi_master_rresp,   --                  .rresp
			h2f_lw_RLAST   => hps_h2f_lw_axi_master_rlast,   --                  .rlast
			h2f_lw_RVALID  => hps_h2f_lw_axi_master_rvalid,  --                  .rvalid
			h2f_lw_RREADY  => hps_h2f_lw_axi_master_rready   --                  .rready
		);

	led_indication_0 : component VideoBox_led_indication_0
		port map (
			clk        => sys_sdram_pll_sys_clk_clk,                             --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,              --               reset.reset_n
			address    => mm_interconnect_2_led_indication_0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_2_led_indication_0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_2_led_indication_0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_2_led_indication_0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_2_led_indication_0_s1_readdata,        --                    .readdata
			out_port   => led_bus_export                                         -- external_connection.export
		);

	sdram_controller : component VideoBox_sdram_controller
		port map (
			clk            => sys_sdram_pll_sys_clk_clk,                                  --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,                   -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_controller_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_controller_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_controller_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_controller_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_controller_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_controller_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_controller_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_controller_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_bus_addr,                                             --  wire.export
			zs_ba          => sdram_bus_ba,                                               --      .export
			zs_cas_n       => sdram_bus_cas_n,                                            --      .export
			zs_cke         => sdram_bus_cke,                                              --      .export
			zs_cs_n        => sdram_bus_cs_n,                                             --      .export
			zs_dq          => sdram_bus_dq,                                               --      .export
			zs_dqm         => sdram_bus_dqm,                                              --      .export
			zs_ras_n       => sdram_bus_ras_n,                                            --      .export
			zs_we_n        => sdram_bus_we_n                                              --      .export
		);

	sys_sdram_pll : component VideoBox_sys_sdram_pll
		port map (
			ref_clk_clk        => ref_clock_clk,                    --      ref_clk.clk
			ref_reset_reset    => hps_h2f_reset_reset_ports_inv,    --    ref_reset.reset
			sys_clk_clk        => sys_sdram_pll_sys_clk_clk,        --      sys_clk.clk
			sdram_clk_clk      => sdram_clock_clk,                  --    sdram_clk.clk
			reset_source_reset => sys_sdram_pll_reset_source_reset  -- reset_source.reset
		);

	vga_pll : component VideoBox_vga_pll
		port map (
			refclk   => sys_sdram_pll_sys_clk_clk,        --  refclk.clk
			rst      => sys_sdram_pll_reset_source_reset, --   reset.reset
			outclk_0 => vga_pll_outclk0_clk,              -- outclk0.clk
			locked   => open                              --  locked.export
		);

	vide_dma_controller : component VideoBox_vide_dma_controller
		port map (
			clk                  => sys_sdram_pll_sys_clk_clk,                                                 --                      clk.clk
			reset                => rst_controller_reset_out_reset,                                            --                    reset.reset
			master_address       => vide_dma_controller_avalon_dma_master_address,                             --        avalon_dma_master.address
			master_waitrequest   => vide_dma_controller_avalon_dma_master_waitrequest,                         --                         .waitrequest
			master_arbiterlock   => vide_dma_controller_avalon_dma_master_lock,                                --                         .lock
			master_read          => vide_dma_controller_avalon_dma_master_read,                                --                         .read
			master_readdata      => vide_dma_controller_avalon_dma_master_readdata,                            --                         .readdata
			master_readdatavalid => vide_dma_controller_avalon_dma_master_readdatavalid,                       --                         .readdatavalid
			slave_address        => mm_interconnect_1_vide_dma_controller_avalon_dma_control_slave_address,    -- avalon_dma_control_slave.address
			slave_byteenable     => mm_interconnect_1_vide_dma_controller_avalon_dma_control_slave_byteenable, --                         .byteenable
			slave_read           => mm_interconnect_1_vide_dma_controller_avalon_dma_control_slave_read,       --                         .read
			slave_write          => mm_interconnect_1_vide_dma_controller_avalon_dma_control_slave_write,      --                         .write
			slave_writedata      => mm_interconnect_1_vide_dma_controller_avalon_dma_control_slave_writedata,  --                         .writedata
			slave_readdata       => mm_interconnect_1_vide_dma_controller_avalon_dma_control_slave_readdata,   --                         .readdata
			stream_ready         => vide_dma_controller_avalon_pixel_source_ready,                             --      avalon_pixel_source.ready
			stream_data          => vide_dma_controller_avalon_pixel_source_data,                              --                         .data
			stream_startofpacket => vide_dma_controller_avalon_pixel_source_startofpacket,                     --                         .startofpacket
			stream_endofpacket   => vide_dma_controller_avalon_pixel_source_endofpacket,                       --                         .endofpacket
			stream_valid         => vide_dma_controller_avalon_pixel_source_valid                              --                         .valid
		);

	vide_dma_controller_citanje : component VideoBox_vide_dma_controller_CITANJE
		port map (
			clk                  => sys_sdram_pll_sys_clk_clk,                                                         --                      clk.clk
			reset                => rst_controller_reset_out_reset,                                                    --                    reset.reset
			master_address       => vide_dma_controller_citanje_avalon_dma_master_address,                             --        avalon_dma_master.address
			master_waitrequest   => vide_dma_controller_citanje_avalon_dma_master_waitrequest,                         --                         .waitrequest
			master_arbiterlock   => vide_dma_controller_citanje_avalon_dma_master_lock,                                --                         .lock
			master_read          => vide_dma_controller_citanje_avalon_dma_master_read,                                --                         .read
			master_readdata      => vide_dma_controller_citanje_avalon_dma_master_readdata,                            --                         .readdata
			master_readdatavalid => vide_dma_controller_citanje_avalon_dma_master_readdatavalid,                       --                         .readdatavalid
			slave_address        => mm_interconnect_1_vide_dma_controller_citanje_avalon_dma_control_slave_address,    -- avalon_dma_control_slave.address
			slave_byteenable     => mm_interconnect_1_vide_dma_controller_citanje_avalon_dma_control_slave_byteenable, --                         .byteenable
			slave_read           => mm_interconnect_1_vide_dma_controller_citanje_avalon_dma_control_slave_read,       --                         .read
			slave_write          => mm_interconnect_1_vide_dma_controller_citanje_avalon_dma_control_slave_write,      --                         .write
			slave_writedata      => mm_interconnect_1_vide_dma_controller_citanje_avalon_dma_control_slave_writedata,  --                         .writedata
			slave_readdata       => mm_interconnect_1_vide_dma_controller_citanje_avalon_dma_control_slave_readdata,   --                         .readdata
			stream_ready         => vide_dma_controller_citanje_avalon_pixel_source_ready,                             --      avalon_pixel_source.ready
			stream_data          => vide_dma_controller_citanje_avalon_pixel_source_data,                              --                         .data
			stream_startofpacket => vide_dma_controller_citanje_avalon_pixel_source_startofpacket,                     --                         .startofpacket
			stream_endofpacket   => vide_dma_controller_citanje_avalon_pixel_source_endofpacket,                       --                         .endofpacket
			stream_valid         => vide_dma_controller_citanje_avalon_pixel_source_valid                              --                         .valid
		);

	vide_dma_controller_citanje_0 : component VideoBox_vide_dma_controller_CITANJE
		port map (
			clk                  => sys_sdram_pll_sys_clk_clk,                                                           --                      clk.clk
			reset                => rst_controller_reset_out_reset,                                                      --                    reset.reset
			master_address       => vide_dma_controller_citanje_0_avalon_dma_master_address,                             --        avalon_dma_master.address
			master_waitrequest   => vide_dma_controller_citanje_0_avalon_dma_master_waitrequest,                         --                         .waitrequest
			master_arbiterlock   => vide_dma_controller_citanje_0_avalon_dma_master_lock,                                --                         .lock
			master_read          => vide_dma_controller_citanje_0_avalon_dma_master_read,                                --                         .read
			master_readdata      => vide_dma_controller_citanje_0_avalon_dma_master_readdata,                            --                         .readdata
			master_readdatavalid => vide_dma_controller_citanje_0_avalon_dma_master_readdatavalid,                       --                         .readdatavalid
			slave_address        => mm_interconnect_1_vide_dma_controller_citanje_0_avalon_dma_control_slave_address,    -- avalon_dma_control_slave.address
			slave_byteenable     => mm_interconnect_1_vide_dma_controller_citanje_0_avalon_dma_control_slave_byteenable, --                         .byteenable
			slave_read           => mm_interconnect_1_vide_dma_controller_citanje_0_avalon_dma_control_slave_read,       --                         .read
			slave_write          => mm_interconnect_1_vide_dma_controller_citanje_0_avalon_dma_control_slave_write,      --                         .write
			slave_writedata      => mm_interconnect_1_vide_dma_controller_citanje_0_avalon_dma_control_slave_writedata,  --                         .writedata
			slave_readdata       => mm_interconnect_1_vide_dma_controller_citanje_0_avalon_dma_control_slave_readdata,   --                         .readdata
			stream_ready         => vide_dma_controller_citanje_0_avalon_pixel_source_ready,                             --      avalon_pixel_source.ready
			stream_data          => vide_dma_controller_citanje_0_avalon_pixel_source_data,                              --                         .data
			stream_startofpacket => vide_dma_controller_citanje_0_avalon_pixel_source_startofpacket,                     --                         .startofpacket
			stream_endofpacket   => vide_dma_controller_citanje_0_avalon_pixel_source_endofpacket,                       --                         .endofpacket
			stream_valid         => vide_dma_controller_citanje_0_avalon_pixel_source_valid                              --                         .valid
		);

	video_dual_clock_buffer : component VideoBox_video_dual_clock_buffer
		port map (
			clk_stream_in            => sys_sdram_pll_sys_clk_clk,                                     --         clock_stream_in.clk
			reset_stream_in          => rst_controller_reset_out_reset,                                --         reset_stream_in.reset
			clk_stream_out           => vga_pll_outclk0_clk,                                           --        clock_stream_out.clk
			reset_stream_out         => rst_controller_001_reset_out_reset,                            --        reset_stream_out.reset
			stream_in_ready          => izbor_prikaza_slike_0_out_ready,                               --   avalon_dc_buffer_sink.ready
			stream_in_startofpacket  => izbor_prikaza_slike_0_out_startofpacket,                       --                        .startofpacket
			stream_in_endofpacket    => izbor_prikaza_slike_0_out_endofpacket,                         --                        .endofpacket
			stream_in_valid          => izbor_prikaza_slike_0_out_valid,                               --                        .valid
			stream_in_data           => izbor_prikaza_slike_0_out_data,                                --                        .data
			stream_out_ready         => video_dual_clock_buffer_avalon_dc_buffer_source_ready,         -- avalon_dc_buffer_source.ready
			stream_out_startofpacket => video_dual_clock_buffer_avalon_dc_buffer_source_startofpacket, --                        .startofpacket
			stream_out_endofpacket   => video_dual_clock_buffer_avalon_dc_buffer_source_endofpacket,   --                        .endofpacket
			stream_out_valid         => video_dual_clock_buffer_avalon_dc_buffer_source_valid,         --                        .valid
			stream_out_data          => video_dual_clock_buffer_avalon_dc_buffer_source_data           --                        .data
		);

	video_rgb_resampler_0 : component VideoBox_video_rgb_resampler_0
		port map (
			clk                      => vga_pll_outclk0_clk,                                           --               clk.clk
			reset                    => rst_controller_001_reset_out_reset,                            --             reset.reset
			stream_in_startofpacket  => video_dual_clock_buffer_avalon_dc_buffer_source_startofpacket, --   avalon_rgb_sink.startofpacket
			stream_in_endofpacket    => video_dual_clock_buffer_avalon_dc_buffer_source_endofpacket,   --                  .endofpacket
			stream_in_valid          => video_dual_clock_buffer_avalon_dc_buffer_source_valid,         --                  .valid
			stream_in_ready          => video_dual_clock_buffer_avalon_dc_buffer_source_ready,         --                  .ready
			stream_in_data           => video_dual_clock_buffer_avalon_dc_buffer_source_data,          --                  .data
			stream_out_ready         => video_rgb_resampler_0_avalon_rgb_source_ready,                 -- avalon_rgb_source.ready
			stream_out_startofpacket => video_rgb_resampler_0_avalon_rgb_source_startofpacket,         --                  .startofpacket
			stream_out_endofpacket   => video_rgb_resampler_0_avalon_rgb_source_endofpacket,           --                  .endofpacket
			stream_out_valid         => video_rgb_resampler_0_avalon_rgb_source_valid,                 --                  .valid
			stream_out_data          => video_rgb_resampler_0_avalon_rgb_source_data                   --                  .data
		);

	video_vga_controller : component VideoBox_video_vga_controller
		port map (
			clk           => vga_pll_outclk0_clk,                                   --                clk.clk
			reset         => rst_controller_001_reset_out_reset,                    --              reset.reset
			data          => video_rgb_resampler_0_avalon_rgb_source_data,          --    avalon_vga_sink.data
			startofpacket => video_rgb_resampler_0_avalon_rgb_source_startofpacket, --                   .startofpacket
			endofpacket   => video_rgb_resampler_0_avalon_rgb_source_endofpacket,   --                   .endofpacket
			valid         => video_rgb_resampler_0_avalon_rgb_source_valid,         --                   .valid
			ready         => video_rgb_resampler_0_avalon_rgb_source_ready,         --                   .ready
			VGA_CLK       => vga_bus_CLK,                                           -- external_interface.export
			VGA_HS        => vga_bus_HS,                                            --                   .export
			VGA_VS        => vga_bus_VS,                                            --                   .export
			VGA_BLANK     => vga_bus_BLANK,                                         --                   .export
			VGA_SYNC      => vga_bus_SYNC,                                          --                   .export
			VGA_R         => vga_bus_R,                                             --                   .export
			VGA_G         => vga_bus_G,                                             --                   .export
			VGA_B         => vga_bus_B                                              --                   .export
		);

	mm_interconnect_0 : component VideoBox_mm_interconnect_0
		port map (
			hps_h2f_axi_master_awid                                        => hps_h2f_axi_master_awid,                                       --                                       hps_h2f_axi_master.awid
			hps_h2f_axi_master_awaddr                                      => hps_h2f_axi_master_awaddr,                                     --                                                         .awaddr
			hps_h2f_axi_master_awlen                                       => hps_h2f_axi_master_awlen,                                      --                                                         .awlen
			hps_h2f_axi_master_awsize                                      => hps_h2f_axi_master_awsize,                                     --                                                         .awsize
			hps_h2f_axi_master_awburst                                     => hps_h2f_axi_master_awburst,                                    --                                                         .awburst
			hps_h2f_axi_master_awlock                                      => hps_h2f_axi_master_awlock,                                     --                                                         .awlock
			hps_h2f_axi_master_awcache                                     => hps_h2f_axi_master_awcache,                                    --                                                         .awcache
			hps_h2f_axi_master_awprot                                      => hps_h2f_axi_master_awprot,                                     --                                                         .awprot
			hps_h2f_axi_master_awvalid                                     => hps_h2f_axi_master_awvalid,                                    --                                                         .awvalid
			hps_h2f_axi_master_awready                                     => hps_h2f_axi_master_awready,                                    --                                                         .awready
			hps_h2f_axi_master_wid                                         => hps_h2f_axi_master_wid,                                        --                                                         .wid
			hps_h2f_axi_master_wdata                                       => hps_h2f_axi_master_wdata,                                      --                                                         .wdata
			hps_h2f_axi_master_wstrb                                       => hps_h2f_axi_master_wstrb,                                      --                                                         .wstrb
			hps_h2f_axi_master_wlast                                       => hps_h2f_axi_master_wlast,                                      --                                                         .wlast
			hps_h2f_axi_master_wvalid                                      => hps_h2f_axi_master_wvalid,                                     --                                                         .wvalid
			hps_h2f_axi_master_wready                                      => hps_h2f_axi_master_wready,                                     --                                                         .wready
			hps_h2f_axi_master_bid                                         => hps_h2f_axi_master_bid,                                        --                                                         .bid
			hps_h2f_axi_master_bresp                                       => hps_h2f_axi_master_bresp,                                      --                                                         .bresp
			hps_h2f_axi_master_bvalid                                      => hps_h2f_axi_master_bvalid,                                     --                                                         .bvalid
			hps_h2f_axi_master_bready                                      => hps_h2f_axi_master_bready,                                     --                                                         .bready
			hps_h2f_axi_master_arid                                        => hps_h2f_axi_master_arid,                                       --                                                         .arid
			hps_h2f_axi_master_araddr                                      => hps_h2f_axi_master_araddr,                                     --                                                         .araddr
			hps_h2f_axi_master_arlen                                       => hps_h2f_axi_master_arlen,                                      --                                                         .arlen
			hps_h2f_axi_master_arsize                                      => hps_h2f_axi_master_arsize,                                     --                                                         .arsize
			hps_h2f_axi_master_arburst                                     => hps_h2f_axi_master_arburst,                                    --                                                         .arburst
			hps_h2f_axi_master_arlock                                      => hps_h2f_axi_master_arlock,                                     --                                                         .arlock
			hps_h2f_axi_master_arcache                                     => hps_h2f_axi_master_arcache,                                    --                                                         .arcache
			hps_h2f_axi_master_arprot                                      => hps_h2f_axi_master_arprot,                                     --                                                         .arprot
			hps_h2f_axi_master_arvalid                                     => hps_h2f_axi_master_arvalid,                                    --                                                         .arvalid
			hps_h2f_axi_master_arready                                     => hps_h2f_axi_master_arready,                                    --                                                         .arready
			hps_h2f_axi_master_rid                                         => hps_h2f_axi_master_rid,                                        --                                                         .rid
			hps_h2f_axi_master_rdata                                       => hps_h2f_axi_master_rdata,                                      --                                                         .rdata
			hps_h2f_axi_master_rresp                                       => hps_h2f_axi_master_rresp,                                      --                                                         .rresp
			hps_h2f_axi_master_rlast                                       => hps_h2f_axi_master_rlast,                                      --                                                         .rlast
			hps_h2f_axi_master_rvalid                                      => hps_h2f_axi_master_rvalid,                                     --                                                         .rvalid
			hps_h2f_axi_master_rready                                      => hps_h2f_axi_master_rready,                                     --                                                         .rready
			sys_sdram_pll_sys_clk_clk                                      => sys_sdram_pll_sys_clk_clk,                                     --                                    sys_sdram_pll_sys_clk.clk
			hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,                            -- hps_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			vide_dma_controller_reset_reset_bridge_in_reset_reset          => rst_controller_reset_out_reset,                                --          vide_dma_controller_reset_reset_bridge_in_reset.reset
			dma_afina_matrica_citanje_avalon_dma_master_address            => dma_afina_matrica_citanje_avalon_dma_master_address,           --              dma_afina_matrica_citanje_avalon_dma_master.address
			dma_afina_matrica_citanje_avalon_dma_master_waitrequest        => dma_afina_matrica_citanje_avalon_dma_master_waitrequest,       --                                                         .waitrequest
			dma_afina_matrica_citanje_avalon_dma_master_read               => dma_afina_matrica_citanje_avalon_dma_master_read,              --                                                         .read
			dma_afina_matrica_citanje_avalon_dma_master_readdata           => dma_afina_matrica_citanje_avalon_dma_master_readdata,          --                                                         .readdata
			dma_afina_matrica_citanje_avalon_dma_master_readdatavalid      => dma_afina_matrica_citanje_avalon_dma_master_readdatavalid,     --                                                         .readdatavalid
			dma_afina_matrica_citanje_avalon_dma_master_lock               => dma_afina_matrica_citanje_avalon_dma_master_lock,              --                                                         .lock
			DMA_CONTROLLER_UPIS_avalon_dma_master_address                  => dma_controller_upis_avalon_dma_master_address,                 --                    DMA_CONTROLLER_UPIS_avalon_dma_master.address
			DMA_CONTROLLER_UPIS_avalon_dma_master_waitrequest              => dma_controller_upis_avalon_dma_master_waitrequest,             --                                                         .waitrequest
			DMA_CONTROLLER_UPIS_avalon_dma_master_write                    => dma_controller_upis_avalon_dma_master_write,                   --                                                         .write
			DMA_CONTROLLER_UPIS_avalon_dma_master_writedata                => dma_controller_upis_avalon_dma_master_writedata,               --                                                         .writedata
			vide_dma_controller_avalon_dma_master_address                  => vide_dma_controller_avalon_dma_master_address,                 --                    vide_dma_controller_avalon_dma_master.address
			vide_dma_controller_avalon_dma_master_waitrequest              => vide_dma_controller_avalon_dma_master_waitrequest,             --                                                         .waitrequest
			vide_dma_controller_avalon_dma_master_read                     => vide_dma_controller_avalon_dma_master_read,                    --                                                         .read
			vide_dma_controller_avalon_dma_master_readdata                 => vide_dma_controller_avalon_dma_master_readdata,                --                                                         .readdata
			vide_dma_controller_avalon_dma_master_readdatavalid            => vide_dma_controller_avalon_dma_master_readdatavalid,           --                                                         .readdatavalid
			vide_dma_controller_avalon_dma_master_lock                     => vide_dma_controller_avalon_dma_master_lock,                    --                                                         .lock
			vide_dma_controller_CITANJE_avalon_dma_master_address          => vide_dma_controller_citanje_avalon_dma_master_address,         --            vide_dma_controller_CITANJE_avalon_dma_master.address
			vide_dma_controller_CITANJE_avalon_dma_master_waitrequest      => vide_dma_controller_citanje_avalon_dma_master_waitrequest,     --                                                         .waitrequest
			vide_dma_controller_CITANJE_avalon_dma_master_read             => vide_dma_controller_citanje_avalon_dma_master_read,            --                                                         .read
			vide_dma_controller_CITANJE_avalon_dma_master_readdata         => vide_dma_controller_citanje_avalon_dma_master_readdata,        --                                                         .readdata
			vide_dma_controller_CITANJE_avalon_dma_master_readdatavalid    => vide_dma_controller_citanje_avalon_dma_master_readdatavalid,   --                                                         .readdatavalid
			vide_dma_controller_CITANJE_avalon_dma_master_lock             => vide_dma_controller_citanje_avalon_dma_master_lock,            --                                                         .lock
			vide_dma_controller_CITANJE_0_avalon_dma_master_address        => vide_dma_controller_citanje_0_avalon_dma_master_address,       --          vide_dma_controller_CITANJE_0_avalon_dma_master.address
			vide_dma_controller_CITANJE_0_avalon_dma_master_waitrequest    => vide_dma_controller_citanje_0_avalon_dma_master_waitrequest,   --                                                         .waitrequest
			vide_dma_controller_CITANJE_0_avalon_dma_master_read           => vide_dma_controller_citanje_0_avalon_dma_master_read,          --                                                         .read
			vide_dma_controller_CITANJE_0_avalon_dma_master_readdata       => vide_dma_controller_citanje_0_avalon_dma_master_readdata,      --                                                         .readdata
			vide_dma_controller_CITANJE_0_avalon_dma_master_readdatavalid  => vide_dma_controller_citanje_0_avalon_dma_master_readdatavalid, --                                                         .readdatavalid
			vide_dma_controller_CITANJE_0_avalon_dma_master_lock           => vide_dma_controller_citanje_0_avalon_dma_master_lock,          --                                                         .lock
			affine_matrix_s1_address                                       => mm_interconnect_0_affine_matrix_s1_address,                    --                                         affine_matrix_s1.address
			affine_matrix_s1_write                                         => mm_interconnect_0_affine_matrix_s1_write,                      --                                                         .write
			affine_matrix_s1_readdata                                      => mm_interconnect_0_affine_matrix_s1_readdata,                   --                                                         .readdata
			affine_matrix_s1_writedata                                     => mm_interconnect_0_affine_matrix_s1_writedata,                  --                                                         .writedata
			affine_matrix_s1_byteenable                                    => mm_interconnect_0_affine_matrix_s1_byteenable,                 --                                                         .byteenable
			affine_matrix_s1_chipselect                                    => mm_interconnect_0_affine_matrix_s1_chipselect,                 --                                                         .chipselect
			affine_matrix_s1_clken                                         => mm_interconnect_0_affine_matrix_s1_clken,                      --                                                         .clken
			sdram_controller_s1_address                                    => mm_interconnect_0_sdram_controller_s1_address,                 --                                      sdram_controller_s1.address
			sdram_controller_s1_write                                      => mm_interconnect_0_sdram_controller_s1_write,                   --                                                         .write
			sdram_controller_s1_read                                       => mm_interconnect_0_sdram_controller_s1_read,                    --                                                         .read
			sdram_controller_s1_readdata                                   => mm_interconnect_0_sdram_controller_s1_readdata,                --                                                         .readdata
			sdram_controller_s1_writedata                                  => mm_interconnect_0_sdram_controller_s1_writedata,               --                                                         .writedata
			sdram_controller_s1_byteenable                                 => mm_interconnect_0_sdram_controller_s1_byteenable,              --                                                         .byteenable
			sdram_controller_s1_readdatavalid                              => mm_interconnect_0_sdram_controller_s1_readdatavalid,           --                                                         .readdatavalid
			sdram_controller_s1_waitrequest                                => mm_interconnect_0_sdram_controller_s1_waitrequest,             --                                                         .waitrequest
			sdram_controller_s1_chipselect                                 => mm_interconnect_0_sdram_controller_s1_chipselect               --                                                         .chipselect
		);

	mm_interconnect_1 : component VideoBox_mm_interconnect_1
		port map (
			hps_h2f_lw_axi_master_awid                                        => hps_h2f_lw_axi_master_awid,                                                          --                                       hps_h2f_lw_axi_master.awid
			hps_h2f_lw_axi_master_awaddr                                      => hps_h2f_lw_axi_master_awaddr,                                                        --                                                            .awaddr
			hps_h2f_lw_axi_master_awlen                                       => hps_h2f_lw_axi_master_awlen,                                                         --                                                            .awlen
			hps_h2f_lw_axi_master_awsize                                      => hps_h2f_lw_axi_master_awsize,                                                        --                                                            .awsize
			hps_h2f_lw_axi_master_awburst                                     => hps_h2f_lw_axi_master_awburst,                                                       --                                                            .awburst
			hps_h2f_lw_axi_master_awlock                                      => hps_h2f_lw_axi_master_awlock,                                                        --                                                            .awlock
			hps_h2f_lw_axi_master_awcache                                     => hps_h2f_lw_axi_master_awcache,                                                       --                                                            .awcache
			hps_h2f_lw_axi_master_awprot                                      => hps_h2f_lw_axi_master_awprot,                                                        --                                                            .awprot
			hps_h2f_lw_axi_master_awvalid                                     => hps_h2f_lw_axi_master_awvalid,                                                       --                                                            .awvalid
			hps_h2f_lw_axi_master_awready                                     => hps_h2f_lw_axi_master_awready,                                                       --                                                            .awready
			hps_h2f_lw_axi_master_wid                                         => hps_h2f_lw_axi_master_wid,                                                           --                                                            .wid
			hps_h2f_lw_axi_master_wdata                                       => hps_h2f_lw_axi_master_wdata,                                                         --                                                            .wdata
			hps_h2f_lw_axi_master_wstrb                                       => hps_h2f_lw_axi_master_wstrb,                                                         --                                                            .wstrb
			hps_h2f_lw_axi_master_wlast                                       => hps_h2f_lw_axi_master_wlast,                                                         --                                                            .wlast
			hps_h2f_lw_axi_master_wvalid                                      => hps_h2f_lw_axi_master_wvalid,                                                        --                                                            .wvalid
			hps_h2f_lw_axi_master_wready                                      => hps_h2f_lw_axi_master_wready,                                                        --                                                            .wready
			hps_h2f_lw_axi_master_bid                                         => hps_h2f_lw_axi_master_bid,                                                           --                                                            .bid
			hps_h2f_lw_axi_master_bresp                                       => hps_h2f_lw_axi_master_bresp,                                                         --                                                            .bresp
			hps_h2f_lw_axi_master_bvalid                                      => hps_h2f_lw_axi_master_bvalid,                                                        --                                                            .bvalid
			hps_h2f_lw_axi_master_bready                                      => hps_h2f_lw_axi_master_bready,                                                        --                                                            .bready
			hps_h2f_lw_axi_master_arid                                        => hps_h2f_lw_axi_master_arid,                                                          --                                                            .arid
			hps_h2f_lw_axi_master_araddr                                      => hps_h2f_lw_axi_master_araddr,                                                        --                                                            .araddr
			hps_h2f_lw_axi_master_arlen                                       => hps_h2f_lw_axi_master_arlen,                                                         --                                                            .arlen
			hps_h2f_lw_axi_master_arsize                                      => hps_h2f_lw_axi_master_arsize,                                                        --                                                            .arsize
			hps_h2f_lw_axi_master_arburst                                     => hps_h2f_lw_axi_master_arburst,                                                       --                                                            .arburst
			hps_h2f_lw_axi_master_arlock                                      => hps_h2f_lw_axi_master_arlock,                                                        --                                                            .arlock
			hps_h2f_lw_axi_master_arcache                                     => hps_h2f_lw_axi_master_arcache,                                                       --                                                            .arcache
			hps_h2f_lw_axi_master_arprot                                      => hps_h2f_lw_axi_master_arprot,                                                        --                                                            .arprot
			hps_h2f_lw_axi_master_arvalid                                     => hps_h2f_lw_axi_master_arvalid,                                                       --                                                            .arvalid
			hps_h2f_lw_axi_master_arready                                     => hps_h2f_lw_axi_master_arready,                                                       --                                                            .arready
			hps_h2f_lw_axi_master_rid                                         => hps_h2f_lw_axi_master_rid,                                                           --                                                            .rid
			hps_h2f_lw_axi_master_rdata                                       => hps_h2f_lw_axi_master_rdata,                                                         --                                                            .rdata
			hps_h2f_lw_axi_master_rresp                                       => hps_h2f_lw_axi_master_rresp,                                                         --                                                            .rresp
			hps_h2f_lw_axi_master_rlast                                       => hps_h2f_lw_axi_master_rlast,                                                         --                                                            .rlast
			hps_h2f_lw_axi_master_rvalid                                      => hps_h2f_lw_axi_master_rvalid,                                                        --                                                            .rvalid
			hps_h2f_lw_axi_master_rready                                      => hps_h2f_lw_axi_master_rready,                                                        --                                                            .rready
			sys_sdram_pll_sys_clk_clk                                         => sys_sdram_pll_sys_clk_clk,                                                           --                                       sys_sdram_pll_sys_clk.clk
			hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,                                                  -- hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			vide_dma_controller_reset_reset_bridge_in_reset_reset             => rst_controller_reset_out_reset,                                                      --             vide_dma_controller_reset_reset_bridge_in_reset.reset
			DMA_CONTROLLER_UPIS_avalon_dma_control_slave_address              => mm_interconnect_1_dma_controller_upis_avalon_dma_control_slave_address,              --                DMA_CONTROLLER_UPIS_avalon_dma_control_slave.address
			DMA_CONTROLLER_UPIS_avalon_dma_control_slave_write                => mm_interconnect_1_dma_controller_upis_avalon_dma_control_slave_write,                --                                                            .write
			DMA_CONTROLLER_UPIS_avalon_dma_control_slave_read                 => mm_interconnect_1_dma_controller_upis_avalon_dma_control_slave_read,                 --                                                            .read
			DMA_CONTROLLER_UPIS_avalon_dma_control_slave_readdata             => mm_interconnect_1_dma_controller_upis_avalon_dma_control_slave_readdata,             --                                                            .readdata
			DMA_CONTROLLER_UPIS_avalon_dma_control_slave_writedata            => mm_interconnect_1_dma_controller_upis_avalon_dma_control_slave_writedata,            --                                                            .writedata
			DMA_CONTROLLER_UPIS_avalon_dma_control_slave_byteenable           => mm_interconnect_1_dma_controller_upis_avalon_dma_control_slave_byteenable,           --                                                            .byteenable
			Image_Processing_0_s0_address                                     => mm_interconnect_1_image_processing_0_s0_address,                                     --                                       Image_Processing_0_s0.address
			Image_Processing_0_s0_write                                       => mm_interconnect_1_image_processing_0_s0_write,                                       --                                                            .write
			Image_Processing_0_s0_read                                        => mm_interconnect_1_image_processing_0_s0_read,                                        --                                                            .read
			Image_Processing_0_s0_readdata                                    => mm_interconnect_1_image_processing_0_s0_readdata,                                    --                                                            .readdata
			Image_Processing_0_s0_writedata                                   => mm_interconnect_1_image_processing_0_s0_writedata,                                   --                                                            .writedata
			Izbor_Prikaza_Slike_0_izbor_slike_address                         => mm_interconnect_1_izbor_prikaza_slike_0_izbor_slike_address,                         --                           Izbor_Prikaza_Slike_0_izbor_slike.address
			Izbor_Prikaza_Slike_0_izbor_slike_write                           => mm_interconnect_1_izbor_prikaza_slike_0_izbor_slike_write,                           --                                                            .write
			Izbor_Prikaza_Slike_0_izbor_slike_read                            => mm_interconnect_1_izbor_prikaza_slike_0_izbor_slike_read,                            --                                                            .read
			Izbor_Prikaza_Slike_0_izbor_slike_readdata                        => mm_interconnect_1_izbor_prikaza_slike_0_izbor_slike_readdata,                        --                                                            .readdata
			Izbor_Prikaza_Slike_0_izbor_slike_writedata                       => mm_interconnect_1_izbor_prikaza_slike_0_izbor_slike_writedata,                       --                                                            .writedata
			vide_dma_controller_avalon_dma_control_slave_address              => mm_interconnect_1_vide_dma_controller_avalon_dma_control_slave_address,              --                vide_dma_controller_avalon_dma_control_slave.address
			vide_dma_controller_avalon_dma_control_slave_write                => mm_interconnect_1_vide_dma_controller_avalon_dma_control_slave_write,                --                                                            .write
			vide_dma_controller_avalon_dma_control_slave_read                 => mm_interconnect_1_vide_dma_controller_avalon_dma_control_slave_read,                 --                                                            .read
			vide_dma_controller_avalon_dma_control_slave_readdata             => mm_interconnect_1_vide_dma_controller_avalon_dma_control_slave_readdata,             --                                                            .readdata
			vide_dma_controller_avalon_dma_control_slave_writedata            => mm_interconnect_1_vide_dma_controller_avalon_dma_control_slave_writedata,            --                                                            .writedata
			vide_dma_controller_avalon_dma_control_slave_byteenable           => mm_interconnect_1_vide_dma_controller_avalon_dma_control_slave_byteenable,           --                                                            .byteenable
			vide_dma_controller_CITANJE_avalon_dma_control_slave_address      => mm_interconnect_1_vide_dma_controller_citanje_avalon_dma_control_slave_address,      --        vide_dma_controller_CITANJE_avalon_dma_control_slave.address
			vide_dma_controller_CITANJE_avalon_dma_control_slave_write        => mm_interconnect_1_vide_dma_controller_citanje_avalon_dma_control_slave_write,        --                                                            .write
			vide_dma_controller_CITANJE_avalon_dma_control_slave_read         => mm_interconnect_1_vide_dma_controller_citanje_avalon_dma_control_slave_read,         --                                                            .read
			vide_dma_controller_CITANJE_avalon_dma_control_slave_readdata     => mm_interconnect_1_vide_dma_controller_citanje_avalon_dma_control_slave_readdata,     --                                                            .readdata
			vide_dma_controller_CITANJE_avalon_dma_control_slave_writedata    => mm_interconnect_1_vide_dma_controller_citanje_avalon_dma_control_slave_writedata,    --                                                            .writedata
			vide_dma_controller_CITANJE_avalon_dma_control_slave_byteenable   => mm_interconnect_1_vide_dma_controller_citanje_avalon_dma_control_slave_byteenable,   --                                                            .byteenable
			vide_dma_controller_CITANJE_0_avalon_dma_control_slave_address    => mm_interconnect_1_vide_dma_controller_citanje_0_avalon_dma_control_slave_address,    --      vide_dma_controller_CITANJE_0_avalon_dma_control_slave.address
			vide_dma_controller_CITANJE_0_avalon_dma_control_slave_write      => mm_interconnect_1_vide_dma_controller_citanje_0_avalon_dma_control_slave_write,      --                                                            .write
			vide_dma_controller_CITANJE_0_avalon_dma_control_slave_read       => mm_interconnect_1_vide_dma_controller_citanje_0_avalon_dma_control_slave_read,       --                                                            .read
			vide_dma_controller_CITANJE_0_avalon_dma_control_slave_readdata   => mm_interconnect_1_vide_dma_controller_citanje_0_avalon_dma_control_slave_readdata,   --                                                            .readdata
			vide_dma_controller_CITANJE_0_avalon_dma_control_slave_writedata  => mm_interconnect_1_vide_dma_controller_citanje_0_avalon_dma_control_slave_writedata,  --                                                            .writedata
			vide_dma_controller_CITANJE_0_avalon_dma_control_slave_byteenable => mm_interconnect_1_vide_dma_controller_citanje_0_avalon_dma_control_slave_byteenable  --                                                            .byteenable
		);

	mm_interconnect_2 : component VideoBox_mm_interconnect_2
		port map (
			sys_sdram_pll_sys_clk_clk                               => sys_sdram_pll_sys_clk_clk,                        --                             sys_sdram_pll_sys_clk.clk
			Izbor_Prikaza_Slike_0_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                   -- Izbor_Prikaza_Slike_0_reset_reset_bridge_in_reset.reset
			Izbor_Prikaza_Slike_0_led_master_waitrequest            => izbor_prikaza_slike_0_led_master_waitrequest,     --                  Izbor_Prikaza_Slike_0_led_master.waitrequest
			Izbor_Prikaza_Slike_0_led_master_write                  => izbor_prikaza_slike_0_led_master_write,           --                                                  .write
			Izbor_Prikaza_Slike_0_led_master_writedata              => izbor_prikaza_slike_0_led_master_writedata,       --                                                  .writedata
			led_indication_0_s1_address                             => mm_interconnect_2_led_indication_0_s1_address,    --                               led_indication_0_s1.address
			led_indication_0_s1_write                               => mm_interconnect_2_led_indication_0_s1_write,      --                                                  .write
			led_indication_0_s1_readdata                            => mm_interconnect_2_led_indication_0_s1_readdata,   --                                                  .readdata
			led_indication_0_s1_writedata                           => mm_interconnect_2_led_indication_0_s1_writedata,  --                                                  .writedata
			led_indication_0_s1_chipselect                          => mm_interconnect_2_led_indication_0_s1_chipselect  --                                                  .chipselect
		);

	rst_controller : component videobox_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => sys_sdram_pll_reset_source_reset,   -- reset_in0.reset
			clk            => sys_sdram_pll_sys_clk_clk,          --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component videobox_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => sys_sdram_pll_reset_source_reset,   -- reset_in0.reset
			clk            => vga_pll_outclk0_clk,                --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component videobox_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => hps_h2f_reset_reset_ports_inv,      -- reset_in0.reset
			clk            => sys_sdram_pll_sys_clk_clk,          --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	hps_h2f_reset_reset_ports_inv <= not hps_h2f_reset_reset;

	mm_interconnect_0_sdram_controller_s1_read_ports_inv <= not mm_interconnect_0_sdram_controller_s1_read;

	mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_controller_s1_byteenable;

	mm_interconnect_0_sdram_controller_s1_write_ports_inv <= not mm_interconnect_0_sdram_controller_s1_write;

	mm_interconnect_2_led_indication_0_s1_write_ports_inv <= not mm_interconnect_2_led_indication_0_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of VideoBox
